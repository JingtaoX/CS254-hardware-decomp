

module top
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  yumi_o,
  v_o,
  ready_i
);

  input [5:0] tag_i;
  output [63:0] v_o;
  output [63:0] v_o1; // added for decompiling
  input [63:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;
  output yumi_o1; // added for decompiling

  bsg_1_to_n_tagged
  wrapper
  (
    .tag_i(tag_i),
    .v_o(v_o),
    .ready_i(ready_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_o(yumi_o)
  );

  bsg_1_to_n_tagged
  wrapper1
  (
    .tag_i(tag_i),
    .v_o(v_o1), // added for decompiling
    .ready_i(ready_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_o(yumi_o1) // added for decompiling
  );
  


endmodule



module bsg_decode_num_out_p64
(
  i,
  o
);

  input [5:0] i;
  output [63:0] o;
  wire [63:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_decode_with_v_num_out_p64
(
  i,
  v_i,
  o
);

  input [5:0] i;
  output [63:0] o;
  input v_i;
  wire [63:0] o,lo;

  bsg_decode_num_out_p64
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[63] = v_i & lo[63];
  assign o[62] = v_i & lo[62];
  assign o[61] = v_i & lo[61];
  assign o[60] = v_i & lo[60];
  assign o[59] = v_i & lo[59];
  assign o[58] = v_i & lo[58];
  assign o[57] = v_i & lo[57];
  assign o[56] = v_i & lo[56];
  assign o[55] = v_i & lo[55];
  assign o[54] = v_i & lo[54];
  assign o[53] = v_i & lo[53];
  assign o[52] = v_i & lo[52];
  assign o[51] = v_i & lo[51];
  assign o[50] = v_i & lo[50];
  assign o[49] = v_i & lo[49];
  assign o[48] = v_i & lo[48];
  assign o[47] = v_i & lo[47];
  assign o[46] = v_i & lo[46];
  assign o[45] = v_i & lo[45];
  assign o[44] = v_i & lo[44];
  assign o[43] = v_i & lo[43];
  assign o[42] = v_i & lo[42];
  assign o[41] = v_i & lo[41];
  assign o[40] = v_i & lo[40];
  assign o[39] = v_i & lo[39];
  assign o[38] = v_i & lo[38];
  assign o[37] = v_i & lo[37];
  assign o[36] = v_i & lo[36];
  assign o[35] = v_i & lo[35];
  assign o[34] = v_i & lo[34];
  assign o[33] = v_i & lo[33];
  assign o[32] = v_i & lo[32];
  assign o[31] = v_i & lo[31];
  assign o[30] = v_i & lo[30];
  assign o[29] = v_i & lo[29];
  assign o[28] = v_i & lo[28];
  assign o[27] = v_i & lo[27];
  assign o[26] = v_i & lo[26];
  assign o[25] = v_i & lo[25];
  assign o[24] = v_i & lo[24];
  assign o[23] = v_i & lo[23];
  assign o[22] = v_i & lo[22];
  assign o[21] = v_i & lo[21];
  assign o[20] = v_i & lo[20];
  assign o[19] = v_i & lo[19];
  assign o[18] = v_i & lo[18];
  assign o[17] = v_i & lo[17];
  assign o[16] = v_i & lo[16];
  assign o[15] = v_i & lo[15];
  assign o[14] = v_i & lo[14];
  assign o[13] = v_i & lo[13];
  assign o[12] = v_i & lo[12];
  assign o[11] = v_i & lo[11];
  assign o[10] = v_i & lo[10];
  assign o[9] = v_i & lo[9];
  assign o[8] = v_i & lo[8];
  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bsg_1_to_n_tagged
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  yumi_o,
  v_o,
  ready_i
);

  input [5:0] tag_i;
  output [63:0] v_o;
  input [63:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;
  wire [63:0] v_o;
  wire yumi_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130;

  bsg_decode_with_v_num_out_p64
  \many.bdv 
  (
    .i(tag_i),
    .v_i(v_i),
    .o(v_o)
  );

  assign N130 = (N66)? ready_i[0] : 
                (N68)? ready_i[1] : 
                (N70)? ready_i[2] : 
                (N72)? ready_i[3] : 
                (N74)? ready_i[4] : 
                (N76)? ready_i[5] : 
                (N78)? ready_i[6] : 
                (N80)? ready_i[7] : 
                (N82)? ready_i[8] : 
                (N84)? ready_i[9] : 
                (N86)? ready_i[10] : 
                (N88)? ready_i[11] : 
                (N90)? ready_i[12] : 
                (N92)? ready_i[13] : 
                (N94)? ready_i[14] : 
                (N96)? ready_i[15] : 
                (N98)? ready_i[16] : 
                (N100)? ready_i[17] : 
                (N102)? ready_i[18] : 
                (N104)? ready_i[19] : 
                (N106)? ready_i[20] : 
                (N108)? ready_i[21] : 
                (N110)? ready_i[22] : 
                (N112)? ready_i[23] : 
                (N114)? ready_i[24] : 
                (N116)? ready_i[25] : 
                (N118)? ready_i[26] : 
                (N120)? ready_i[27] : 
                (N122)? ready_i[28] : 
                (N124)? ready_i[29] : 
                (N126)? ready_i[30] : 
                (N128)? ready_i[31] : 
                (N67)? ready_i[32] : 
                (N69)? ready_i[33] : 
                (N71)? ready_i[34] : 
                (N73)? ready_i[35] : 
                (N75)? ready_i[36] : 
                (N77)? ready_i[37] : 
                (N79)? ready_i[38] : 
                (N81)? ready_i[39] : 
                (N83)? ready_i[40] : 
                (N85)? ready_i[41] : 
                (N87)? ready_i[42] : 
                (N89)? ready_i[43] : 
                (N91)? ready_i[44] : 
                (N93)? ready_i[45] : 
                (N95)? ready_i[46] : 
                (N97)? ready_i[47] : 
                (N99)? ready_i[48] : 
                (N101)? ready_i[49] : 
                (N103)? ready_i[50] : 
                (N105)? ready_i[51] : 
                (N107)? ready_i[52] : 
                (N109)? ready_i[53] : 
                (N111)? ready_i[54] : 
                (N113)? ready_i[55] : 
                (N115)? ready_i[56] : 
                (N117)? ready_i[57] : 
                (N119)? ready_i[58] : 
                (N121)? ready_i[59] : 
                (N123)? ready_i[60] : 
                (N125)? ready_i[61] : 
                (N127)? ready_i[62] : 
                (N129)? ready_i[63] : 1'b0;
  assign N0 = ~tag_i[0];
  assign N1 = ~tag_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & tag_i[1];
  assign N4 = tag_i[0] & N1;
  assign N5 = tag_i[0] & tag_i[1];
  assign N6 = ~tag_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & tag_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & tag_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & tag_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & tag_i[2];
  assign N15 = ~tag_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & tag_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & tag_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & tag_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & tag_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & tag_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & tag_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & tag_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & tag_i[3];
  assign N32 = ~tag_i[4];
  assign N33 = N16 & N32;
  assign N34 = N16 & tag_i[4];
  assign N35 = N18 & N32;
  assign N36 = N18 & tag_i[4];
  assign N37 = N20 & N32;
  assign N38 = N20 & tag_i[4];
  assign N39 = N22 & N32;
  assign N40 = N22 & tag_i[4];
  assign N41 = N24 & N32;
  assign N42 = N24 & tag_i[4];
  assign N43 = N26 & N32;
  assign N44 = N26 & tag_i[4];
  assign N45 = N28 & N32;
  assign N46 = N28 & tag_i[4];
  assign N47 = N30 & N32;
  assign N48 = N30 & tag_i[4];
  assign N49 = N17 & N32;
  assign N50 = N17 & tag_i[4];
  assign N51 = N19 & N32;
  assign N52 = N19 & tag_i[4];
  assign N53 = N21 & N32;
  assign N54 = N21 & tag_i[4];
  assign N55 = N23 & N32;
  assign N56 = N23 & tag_i[4];
  assign N57 = N25 & N32;
  assign N58 = N25 & tag_i[4];
  assign N59 = N27 & N32;
  assign N60 = N27 & tag_i[4];
  assign N61 = N29 & N32;
  assign N62 = N29 & tag_i[4];
  assign N63 = N31 & N32;
  assign N64 = N31 & tag_i[4];
  assign N65 = ~tag_i[5];
  assign N66 = N33 & N65;
  assign N67 = N33 & tag_i[5];
  assign N68 = N35 & N65;
  assign N69 = N35 & tag_i[5];
  assign N70 = N37 & N65;
  assign N71 = N37 & tag_i[5];
  assign N72 = N39 & N65;
  assign N73 = N39 & tag_i[5];
  assign N74 = N41 & N65;
  assign N75 = N41 & tag_i[5];
  assign N76 = N43 & N65;
  assign N77 = N43 & tag_i[5];
  assign N78 = N45 & N65;
  assign N79 = N45 & tag_i[5];
  assign N80 = N47 & N65;
  assign N81 = N47 & tag_i[5];
  assign N82 = N49 & N65;
  assign N83 = N49 & tag_i[5];
  assign N84 = N51 & N65;
  assign N85 = N51 & tag_i[5];
  assign N86 = N53 & N65;
  assign N87 = N53 & tag_i[5];
  assign N88 = N55 & N65;
  assign N89 = N55 & tag_i[5];
  assign N90 = N57 & N65;
  assign N91 = N57 & tag_i[5];
  assign N92 = N59 & N65;
  assign N93 = N59 & tag_i[5];
  assign N94 = N61 & N65;
  assign N95 = N61 & tag_i[5];
  assign N96 = N63 & N65;
  assign N97 = N63 & tag_i[5];
  assign N98 = N34 & N65;
  assign N99 = N34 & tag_i[5];
  assign N100 = N36 & N65;
  assign N101 = N36 & tag_i[5];
  assign N102 = N38 & N65;
  assign N103 = N38 & tag_i[5];
  assign N104 = N40 & N65;
  assign N105 = N40 & tag_i[5];
  assign N106 = N42 & N65;
  assign N107 = N42 & tag_i[5];
  assign N108 = N44 & N65;
  assign N109 = N44 & tag_i[5];
  assign N110 = N46 & N65;
  assign N111 = N46 & tag_i[5];
  assign N112 = N48 & N65;
  assign N113 = N48 & tag_i[5];
  assign N114 = N50 & N65;
  assign N115 = N50 & tag_i[5];
  assign N116 = N52 & N65;
  assign N117 = N52 & tag_i[5];
  assign N118 = N54 & N65;
  assign N119 = N54 & tag_i[5];
  assign N120 = N56 & N65;
  assign N121 = N56 & tag_i[5];
  assign N122 = N58 & N65;
  assign N123 = N58 & tag_i[5];
  assign N124 = N60 & N65;
  assign N125 = N60 & tag_i[5];
  assign N126 = N62 & N65;
  assign N127 = N62 & tag_i[5];
  assign N128 = N64 & N65;
  assign N129 = N64 & tag_i[5];
  assign yumi_o = N130 & v_i;

endmodule

