

module top
(
  data_i,
  sel_i,
  data_o,
  data_o1 // added for decompiling
);

  input [511:0] data_i;
  input [4:0] sel_i;
  output [511:0] data_o;
  output [511:0] data_o1; // added for decompiling

  bsg_mux_butterfly
  wrapper
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o)
  );

  bsg_mux_butterfly
  wrapper1
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o1) // added for decompiling
  );


endmodule



module bsg_swap_width_p16
(
  data_i,
  swap_i,
  data_o
);

  input [31:0] data_i;
  output [31:0] data_o;
  input swap_i;
  wire [31:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[15:0], data_i[31:16] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p32
(
  data_i,
  swap_i,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input swap_i;
  wire [63:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[31:0], data_i[63:32] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p64
(
  data_i,
  swap_i,
  data_o
);

  input [127:0] data_i;
  output [127:0] data_o;
  input swap_i;
  wire [127:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[63:0], data_i[127:64] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p128
(
  data_i,
  swap_i,
  data_o
);

  input [255:0] data_i;
  output [255:0] data_o;
  input swap_i;
  wire [255:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[127:0], data_i[255:128] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p256
(
  data_i,
  swap_i,
  data_o
);

  input [511:0] data_i;
  output [511:0] data_o;
  input swap_i;
  wire [511:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[255:0], data_i[511:256] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_mux_butterfly
(
  data_i,
  sel_i,
  data_o
);

  input [511:0] data_i;
  input [4:0] sel_i;
  output [511:0] data_o;
  wire [511:0] data_o;
  wire data_stage_1__511_,data_stage_1__510_,data_stage_1__509_,data_stage_1__508_,
  data_stage_1__507_,data_stage_1__506_,data_stage_1__505_,data_stage_1__504_,
  data_stage_1__503_,data_stage_1__502_,data_stage_1__501_,data_stage_1__500_,
  data_stage_1__499_,data_stage_1__498_,data_stage_1__497_,data_stage_1__496_,
  data_stage_1__495_,data_stage_1__494_,data_stage_1__493_,data_stage_1__492_,data_stage_1__491_,
  data_stage_1__490_,data_stage_1__489_,data_stage_1__488_,data_stage_1__487_,
  data_stage_1__486_,data_stage_1__485_,data_stage_1__484_,data_stage_1__483_,
  data_stage_1__482_,data_stage_1__481_,data_stage_1__480_,data_stage_1__479_,
  data_stage_1__478_,data_stage_1__477_,data_stage_1__476_,data_stage_1__475_,
  data_stage_1__474_,data_stage_1__473_,data_stage_1__472_,data_stage_1__471_,data_stage_1__470_,
  data_stage_1__469_,data_stage_1__468_,data_stage_1__467_,data_stage_1__466_,
  data_stage_1__465_,data_stage_1__464_,data_stage_1__463_,data_stage_1__462_,
  data_stage_1__461_,data_stage_1__460_,data_stage_1__459_,data_stage_1__458_,
  data_stage_1__457_,data_stage_1__456_,data_stage_1__455_,data_stage_1__454_,
  data_stage_1__453_,data_stage_1__452_,data_stage_1__451_,data_stage_1__450_,data_stage_1__449_,
  data_stage_1__448_,data_stage_1__447_,data_stage_1__446_,data_stage_1__445_,
  data_stage_1__444_,data_stage_1__443_,data_stage_1__442_,data_stage_1__441_,
  data_stage_1__440_,data_stage_1__439_,data_stage_1__438_,data_stage_1__437_,
  data_stage_1__436_,data_stage_1__435_,data_stage_1__434_,data_stage_1__433_,data_stage_1__432_,
  data_stage_1__431_,data_stage_1__430_,data_stage_1__429_,data_stage_1__428_,
  data_stage_1__427_,data_stage_1__426_,data_stage_1__425_,data_stage_1__424_,
  data_stage_1__423_,data_stage_1__422_,data_stage_1__421_,data_stage_1__420_,
  data_stage_1__419_,data_stage_1__418_,data_stage_1__417_,data_stage_1__416_,
  data_stage_1__415_,data_stage_1__414_,data_stage_1__413_,data_stage_1__412_,data_stage_1__411_,
  data_stage_1__410_,data_stage_1__409_,data_stage_1__408_,data_stage_1__407_,
  data_stage_1__406_,data_stage_1__405_,data_stage_1__404_,data_stage_1__403_,
  data_stage_1__402_,data_stage_1__401_,data_stage_1__400_,data_stage_1__399_,
  data_stage_1__398_,data_stage_1__397_,data_stage_1__396_,data_stage_1__395_,
  data_stage_1__394_,data_stage_1__393_,data_stage_1__392_,data_stage_1__391_,data_stage_1__390_,
  data_stage_1__389_,data_stage_1__388_,data_stage_1__387_,data_stage_1__386_,
  data_stage_1__385_,data_stage_1__384_,data_stage_1__383_,data_stage_1__382_,
  data_stage_1__381_,data_stage_1__380_,data_stage_1__379_,data_stage_1__378_,
  data_stage_1__377_,data_stage_1__376_,data_stage_1__375_,data_stage_1__374_,
  data_stage_1__373_,data_stage_1__372_,data_stage_1__371_,data_stage_1__370_,data_stage_1__369_,
  data_stage_1__368_,data_stage_1__367_,data_stage_1__366_,data_stage_1__365_,
  data_stage_1__364_,data_stage_1__363_,data_stage_1__362_,data_stage_1__361_,
  data_stage_1__360_,data_stage_1__359_,data_stage_1__358_,data_stage_1__357_,
  data_stage_1__356_,data_stage_1__355_,data_stage_1__354_,data_stage_1__353_,data_stage_1__352_,
  data_stage_1__351_,data_stage_1__350_,data_stage_1__349_,data_stage_1__348_,
  data_stage_1__347_,data_stage_1__346_,data_stage_1__345_,data_stage_1__344_,
  data_stage_1__343_,data_stage_1__342_,data_stage_1__341_,data_stage_1__340_,
  data_stage_1__339_,data_stage_1__338_,data_stage_1__337_,data_stage_1__336_,
  data_stage_1__335_,data_stage_1__334_,data_stage_1__333_,data_stage_1__332_,data_stage_1__331_,
  data_stage_1__330_,data_stage_1__329_,data_stage_1__328_,data_stage_1__327_,
  data_stage_1__326_,data_stage_1__325_,data_stage_1__324_,data_stage_1__323_,
  data_stage_1__322_,data_stage_1__321_,data_stage_1__320_,data_stage_1__319_,
  data_stage_1__318_,data_stage_1__317_,data_stage_1__316_,data_stage_1__315_,
  data_stage_1__314_,data_stage_1__313_,data_stage_1__312_,data_stage_1__311_,data_stage_1__310_,
  data_stage_1__309_,data_stage_1__308_,data_stage_1__307_,data_stage_1__306_,
  data_stage_1__305_,data_stage_1__304_,data_stage_1__303_,data_stage_1__302_,
  data_stage_1__301_,data_stage_1__300_,data_stage_1__299_,data_stage_1__298_,
  data_stage_1__297_,data_stage_1__296_,data_stage_1__295_,data_stage_1__294_,
  data_stage_1__293_,data_stage_1__292_,data_stage_1__291_,data_stage_1__290_,data_stage_1__289_,
  data_stage_1__288_,data_stage_1__287_,data_stage_1__286_,data_stage_1__285_,
  data_stage_1__284_,data_stage_1__283_,data_stage_1__282_,data_stage_1__281_,
  data_stage_1__280_,data_stage_1__279_,data_stage_1__278_,data_stage_1__277_,
  data_stage_1__276_,data_stage_1__275_,data_stage_1__274_,data_stage_1__273_,data_stage_1__272_,
  data_stage_1__271_,data_stage_1__270_,data_stage_1__269_,data_stage_1__268_,
  data_stage_1__267_,data_stage_1__266_,data_stage_1__265_,data_stage_1__264_,
  data_stage_1__263_,data_stage_1__262_,data_stage_1__261_,data_stage_1__260_,
  data_stage_1__259_,data_stage_1__258_,data_stage_1__257_,data_stage_1__256_,
  data_stage_1__255_,data_stage_1__254_,data_stage_1__253_,data_stage_1__252_,data_stage_1__251_,
  data_stage_1__250_,data_stage_1__249_,data_stage_1__248_,data_stage_1__247_,
  data_stage_1__246_,data_stage_1__245_,data_stage_1__244_,data_stage_1__243_,
  data_stage_1__242_,data_stage_1__241_,data_stage_1__240_,data_stage_1__239_,
  data_stage_1__238_,data_stage_1__237_,data_stage_1__236_,data_stage_1__235_,
  data_stage_1__234_,data_stage_1__233_,data_stage_1__232_,data_stage_1__231_,data_stage_1__230_,
  data_stage_1__229_,data_stage_1__228_,data_stage_1__227_,data_stage_1__226_,
  data_stage_1__225_,data_stage_1__224_,data_stage_1__223_,data_stage_1__222_,
  data_stage_1__221_,data_stage_1__220_,data_stage_1__219_,data_stage_1__218_,
  data_stage_1__217_,data_stage_1__216_,data_stage_1__215_,data_stage_1__214_,
  data_stage_1__213_,data_stage_1__212_,data_stage_1__211_,data_stage_1__210_,data_stage_1__209_,
  data_stage_1__208_,data_stage_1__207_,data_stage_1__206_,data_stage_1__205_,
  data_stage_1__204_,data_stage_1__203_,data_stage_1__202_,data_stage_1__201_,
  data_stage_1__200_,data_stage_1__199_,data_stage_1__198_,data_stage_1__197_,
  data_stage_1__196_,data_stage_1__195_,data_stage_1__194_,data_stage_1__193_,data_stage_1__192_,
  data_stage_1__191_,data_stage_1__190_,data_stage_1__189_,data_stage_1__188_,
  data_stage_1__187_,data_stage_1__186_,data_stage_1__185_,data_stage_1__184_,
  data_stage_1__183_,data_stage_1__182_,data_stage_1__181_,data_stage_1__180_,
  data_stage_1__179_,data_stage_1__178_,data_stage_1__177_,data_stage_1__176_,
  data_stage_1__175_,data_stage_1__174_,data_stage_1__173_,data_stage_1__172_,data_stage_1__171_,
  data_stage_1__170_,data_stage_1__169_,data_stage_1__168_,data_stage_1__167_,
  data_stage_1__166_,data_stage_1__165_,data_stage_1__164_,data_stage_1__163_,
  data_stage_1__162_,data_stage_1__161_,data_stage_1__160_,data_stage_1__159_,
  data_stage_1__158_,data_stage_1__157_,data_stage_1__156_,data_stage_1__155_,
  data_stage_1__154_,data_stage_1__153_,data_stage_1__152_,data_stage_1__151_,data_stage_1__150_,
  data_stage_1__149_,data_stage_1__148_,data_stage_1__147_,data_stage_1__146_,
  data_stage_1__145_,data_stage_1__144_,data_stage_1__143_,data_stage_1__142_,
  data_stage_1__141_,data_stage_1__140_,data_stage_1__139_,data_stage_1__138_,
  data_stage_1__137_,data_stage_1__136_,data_stage_1__135_,data_stage_1__134_,
  data_stage_1__133_,data_stage_1__132_,data_stage_1__131_,data_stage_1__130_,data_stage_1__129_,
  data_stage_1__128_,data_stage_1__127_,data_stage_1__126_,data_stage_1__125_,
  data_stage_1__124_,data_stage_1__123_,data_stage_1__122_,data_stage_1__121_,
  data_stage_1__120_,data_stage_1__119_,data_stage_1__118_,data_stage_1__117_,
  data_stage_1__116_,data_stage_1__115_,data_stage_1__114_,data_stage_1__113_,data_stage_1__112_,
  data_stage_1__111_,data_stage_1__110_,data_stage_1__109_,data_stage_1__108_,
  data_stage_1__107_,data_stage_1__106_,data_stage_1__105_,data_stage_1__104_,
  data_stage_1__103_,data_stage_1__102_,data_stage_1__101_,data_stage_1__100_,
  data_stage_1__99_,data_stage_1__98_,data_stage_1__97_,data_stage_1__96_,data_stage_1__95_,
  data_stage_1__94_,data_stage_1__93_,data_stage_1__92_,data_stage_1__91_,
  data_stage_1__90_,data_stage_1__89_,data_stage_1__88_,data_stage_1__87_,data_stage_1__86_,
  data_stage_1__85_,data_stage_1__84_,data_stage_1__83_,data_stage_1__82_,
  data_stage_1__81_,data_stage_1__80_,data_stage_1__79_,data_stage_1__78_,
  data_stage_1__77_,data_stage_1__76_,data_stage_1__75_,data_stage_1__74_,data_stage_1__73_,
  data_stage_1__72_,data_stage_1__71_,data_stage_1__70_,data_stage_1__69_,
  data_stage_1__68_,data_stage_1__67_,data_stage_1__66_,data_stage_1__65_,data_stage_1__64_,
  data_stage_1__63_,data_stage_1__62_,data_stage_1__61_,data_stage_1__60_,
  data_stage_1__59_,data_stage_1__58_,data_stage_1__57_,data_stage_1__56_,data_stage_1__55_,
  data_stage_1__54_,data_stage_1__53_,data_stage_1__52_,data_stage_1__51_,
  data_stage_1__50_,data_stage_1__49_,data_stage_1__48_,data_stage_1__47_,data_stage_1__46_,
  data_stage_1__45_,data_stage_1__44_,data_stage_1__43_,data_stage_1__42_,
  data_stage_1__41_,data_stage_1__40_,data_stage_1__39_,data_stage_1__38_,
  data_stage_1__37_,data_stage_1__36_,data_stage_1__35_,data_stage_1__34_,data_stage_1__33_,
  data_stage_1__32_,data_stage_1__31_,data_stage_1__30_,data_stage_1__29_,
  data_stage_1__28_,data_stage_1__27_,data_stage_1__26_,data_stage_1__25_,data_stage_1__24_,
  data_stage_1__23_,data_stage_1__22_,data_stage_1__21_,data_stage_1__20_,
  data_stage_1__19_,data_stage_1__18_,data_stage_1__17_,data_stage_1__16_,data_stage_1__15_,
  data_stage_1__14_,data_stage_1__13_,data_stage_1__12_,data_stage_1__11_,
  data_stage_1__10_,data_stage_1__9_,data_stage_1__8_,data_stage_1__7_,data_stage_1__6_,
  data_stage_1__5_,data_stage_1__4_,data_stage_1__3_,data_stage_1__2_,
  data_stage_1__1_,data_stage_1__0_,data_stage_2__511_,data_stage_2__510_,data_stage_2__509_,
  data_stage_2__508_,data_stage_2__507_,data_stage_2__506_,data_stage_2__505_,
  data_stage_2__504_,data_stage_2__503_,data_stage_2__502_,data_stage_2__501_,
  data_stage_2__500_,data_stage_2__499_,data_stage_2__498_,data_stage_2__497_,
  data_stage_2__496_,data_stage_2__495_,data_stage_2__494_,data_stage_2__493_,data_stage_2__492_,
  data_stage_2__491_,data_stage_2__490_,data_stage_2__489_,data_stage_2__488_,
  data_stage_2__487_,data_stage_2__486_,data_stage_2__485_,data_stage_2__484_,
  data_stage_2__483_,data_stage_2__482_,data_stage_2__481_,data_stage_2__480_,
  data_stage_2__479_,data_stage_2__478_,data_stage_2__477_,data_stage_2__476_,
  data_stage_2__475_,data_stage_2__474_,data_stage_2__473_,data_stage_2__472_,data_stage_2__471_,
  data_stage_2__470_,data_stage_2__469_,data_stage_2__468_,data_stage_2__467_,
  data_stage_2__466_,data_stage_2__465_,data_stage_2__464_,data_stage_2__463_,
  data_stage_2__462_,data_stage_2__461_,data_stage_2__460_,data_stage_2__459_,
  data_stage_2__458_,data_stage_2__457_,data_stage_2__456_,data_stage_2__455_,data_stage_2__454_,
  data_stage_2__453_,data_stage_2__452_,data_stage_2__451_,data_stage_2__450_,
  data_stage_2__449_,data_stage_2__448_,data_stage_2__447_,data_stage_2__446_,
  data_stage_2__445_,data_stage_2__444_,data_stage_2__443_,data_stage_2__442_,
  data_stage_2__441_,data_stage_2__440_,data_stage_2__439_,data_stage_2__438_,
  data_stage_2__437_,data_stage_2__436_,data_stage_2__435_,data_stage_2__434_,data_stage_2__433_,
  data_stage_2__432_,data_stage_2__431_,data_stage_2__430_,data_stage_2__429_,
  data_stage_2__428_,data_stage_2__427_,data_stage_2__426_,data_stage_2__425_,
  data_stage_2__424_,data_stage_2__423_,data_stage_2__422_,data_stage_2__421_,
  data_stage_2__420_,data_stage_2__419_,data_stage_2__418_,data_stage_2__417_,
  data_stage_2__416_,data_stage_2__415_,data_stage_2__414_,data_stage_2__413_,data_stage_2__412_,
  data_stage_2__411_,data_stage_2__410_,data_stage_2__409_,data_stage_2__408_,
  data_stage_2__407_,data_stage_2__406_,data_stage_2__405_,data_stage_2__404_,
  data_stage_2__403_,data_stage_2__402_,data_stage_2__401_,data_stage_2__400_,
  data_stage_2__399_,data_stage_2__398_,data_stage_2__397_,data_stage_2__396_,
  data_stage_2__395_,data_stage_2__394_,data_stage_2__393_,data_stage_2__392_,data_stage_2__391_,
  data_stage_2__390_,data_stage_2__389_,data_stage_2__388_,data_stage_2__387_,
  data_stage_2__386_,data_stage_2__385_,data_stage_2__384_,data_stage_2__383_,
  data_stage_2__382_,data_stage_2__381_,data_stage_2__380_,data_stage_2__379_,
  data_stage_2__378_,data_stage_2__377_,data_stage_2__376_,data_stage_2__375_,data_stage_2__374_,
  data_stage_2__373_,data_stage_2__372_,data_stage_2__371_,data_stage_2__370_,
  data_stage_2__369_,data_stage_2__368_,data_stage_2__367_,data_stage_2__366_,
  data_stage_2__365_,data_stage_2__364_,data_stage_2__363_,data_stage_2__362_,
  data_stage_2__361_,data_stage_2__360_,data_stage_2__359_,data_stage_2__358_,
  data_stage_2__357_,data_stage_2__356_,data_stage_2__355_,data_stage_2__354_,data_stage_2__353_,
  data_stage_2__352_,data_stage_2__351_,data_stage_2__350_,data_stage_2__349_,
  data_stage_2__348_,data_stage_2__347_,data_stage_2__346_,data_stage_2__345_,
  data_stage_2__344_,data_stage_2__343_,data_stage_2__342_,data_stage_2__341_,
  data_stage_2__340_,data_stage_2__339_,data_stage_2__338_,data_stage_2__337_,
  data_stage_2__336_,data_stage_2__335_,data_stage_2__334_,data_stage_2__333_,data_stage_2__332_,
  data_stage_2__331_,data_stage_2__330_,data_stage_2__329_,data_stage_2__328_,
  data_stage_2__327_,data_stage_2__326_,data_stage_2__325_,data_stage_2__324_,
  data_stage_2__323_,data_stage_2__322_,data_stage_2__321_,data_stage_2__320_,
  data_stage_2__319_,data_stage_2__318_,data_stage_2__317_,data_stage_2__316_,
  data_stage_2__315_,data_stage_2__314_,data_stage_2__313_,data_stage_2__312_,data_stage_2__311_,
  data_stage_2__310_,data_stage_2__309_,data_stage_2__308_,data_stage_2__307_,
  data_stage_2__306_,data_stage_2__305_,data_stage_2__304_,data_stage_2__303_,
  data_stage_2__302_,data_stage_2__301_,data_stage_2__300_,data_stage_2__299_,
  data_stage_2__298_,data_stage_2__297_,data_stage_2__296_,data_stage_2__295_,data_stage_2__294_,
  data_stage_2__293_,data_stage_2__292_,data_stage_2__291_,data_stage_2__290_,
  data_stage_2__289_,data_stage_2__288_,data_stage_2__287_,data_stage_2__286_,
  data_stage_2__285_,data_stage_2__284_,data_stage_2__283_,data_stage_2__282_,
  data_stage_2__281_,data_stage_2__280_,data_stage_2__279_,data_stage_2__278_,
  data_stage_2__277_,data_stage_2__276_,data_stage_2__275_,data_stage_2__274_,data_stage_2__273_,
  data_stage_2__272_,data_stage_2__271_,data_stage_2__270_,data_stage_2__269_,
  data_stage_2__268_,data_stage_2__267_,data_stage_2__266_,data_stage_2__265_,
  data_stage_2__264_,data_stage_2__263_,data_stage_2__262_,data_stage_2__261_,
  data_stage_2__260_,data_stage_2__259_,data_stage_2__258_,data_stage_2__257_,
  data_stage_2__256_,data_stage_2__255_,data_stage_2__254_,data_stage_2__253_,data_stage_2__252_,
  data_stage_2__251_,data_stage_2__250_,data_stage_2__249_,data_stage_2__248_,
  data_stage_2__247_,data_stage_2__246_,data_stage_2__245_,data_stage_2__244_,
  data_stage_2__243_,data_stage_2__242_,data_stage_2__241_,data_stage_2__240_,
  data_stage_2__239_,data_stage_2__238_,data_stage_2__237_,data_stage_2__236_,
  data_stage_2__235_,data_stage_2__234_,data_stage_2__233_,data_stage_2__232_,data_stage_2__231_,
  data_stage_2__230_,data_stage_2__229_,data_stage_2__228_,data_stage_2__227_,
  data_stage_2__226_,data_stage_2__225_,data_stage_2__224_,data_stage_2__223_,
  data_stage_2__222_,data_stage_2__221_,data_stage_2__220_,data_stage_2__219_,
  data_stage_2__218_,data_stage_2__217_,data_stage_2__216_,data_stage_2__215_,data_stage_2__214_,
  data_stage_2__213_,data_stage_2__212_,data_stage_2__211_,data_stage_2__210_,
  data_stage_2__209_,data_stage_2__208_,data_stage_2__207_,data_stage_2__206_,
  data_stage_2__205_,data_stage_2__204_,data_stage_2__203_,data_stage_2__202_,
  data_stage_2__201_,data_stage_2__200_,data_stage_2__199_,data_stage_2__198_,
  data_stage_2__197_,data_stage_2__196_,data_stage_2__195_,data_stage_2__194_,data_stage_2__193_,
  data_stage_2__192_,data_stage_2__191_,data_stage_2__190_,data_stage_2__189_,
  data_stage_2__188_,data_stage_2__187_,data_stage_2__186_,data_stage_2__185_,
  data_stage_2__184_,data_stage_2__183_,data_stage_2__182_,data_stage_2__181_,
  data_stage_2__180_,data_stage_2__179_,data_stage_2__178_,data_stage_2__177_,
  data_stage_2__176_,data_stage_2__175_,data_stage_2__174_,data_stage_2__173_,data_stage_2__172_,
  data_stage_2__171_,data_stage_2__170_,data_stage_2__169_,data_stage_2__168_,
  data_stage_2__167_,data_stage_2__166_,data_stage_2__165_,data_stage_2__164_,
  data_stage_2__163_,data_stage_2__162_,data_stage_2__161_,data_stage_2__160_,
  data_stage_2__159_,data_stage_2__158_,data_stage_2__157_,data_stage_2__156_,
  data_stage_2__155_,data_stage_2__154_,data_stage_2__153_,data_stage_2__152_,data_stage_2__151_,
  data_stage_2__150_,data_stage_2__149_,data_stage_2__148_,data_stage_2__147_,
  data_stage_2__146_,data_stage_2__145_,data_stage_2__144_,data_stage_2__143_,
  data_stage_2__142_,data_stage_2__141_,data_stage_2__140_,data_stage_2__139_,
  data_stage_2__138_,data_stage_2__137_,data_stage_2__136_,data_stage_2__135_,data_stage_2__134_,
  data_stage_2__133_,data_stage_2__132_,data_stage_2__131_,data_stage_2__130_,
  data_stage_2__129_,data_stage_2__128_,data_stage_2__127_,data_stage_2__126_,
  data_stage_2__125_,data_stage_2__124_,data_stage_2__123_,data_stage_2__122_,
  data_stage_2__121_,data_stage_2__120_,data_stage_2__119_,data_stage_2__118_,
  data_stage_2__117_,data_stage_2__116_,data_stage_2__115_,data_stage_2__114_,data_stage_2__113_,
  data_stage_2__112_,data_stage_2__111_,data_stage_2__110_,data_stage_2__109_,
  data_stage_2__108_,data_stage_2__107_,data_stage_2__106_,data_stage_2__105_,
  data_stage_2__104_,data_stage_2__103_,data_stage_2__102_,data_stage_2__101_,
  data_stage_2__100_,data_stage_2__99_,data_stage_2__98_,data_stage_2__97_,data_stage_2__96_,
  data_stage_2__95_,data_stage_2__94_,data_stage_2__93_,data_stage_2__92_,
  data_stage_2__91_,data_stage_2__90_,data_stage_2__89_,data_stage_2__88_,data_stage_2__87_,
  data_stage_2__86_,data_stage_2__85_,data_stage_2__84_,data_stage_2__83_,
  data_stage_2__82_,data_stage_2__81_,data_stage_2__80_,data_stage_2__79_,
  data_stage_2__78_,data_stage_2__77_,data_stage_2__76_,data_stage_2__75_,data_stage_2__74_,
  data_stage_2__73_,data_stage_2__72_,data_stage_2__71_,data_stage_2__70_,
  data_stage_2__69_,data_stage_2__68_,data_stage_2__67_,data_stage_2__66_,data_stage_2__65_,
  data_stage_2__64_,data_stage_2__63_,data_stage_2__62_,data_stage_2__61_,
  data_stage_2__60_,data_stage_2__59_,data_stage_2__58_,data_stage_2__57_,data_stage_2__56_,
  data_stage_2__55_,data_stage_2__54_,data_stage_2__53_,data_stage_2__52_,
  data_stage_2__51_,data_stage_2__50_,data_stage_2__49_,data_stage_2__48_,data_stage_2__47_,
  data_stage_2__46_,data_stage_2__45_,data_stage_2__44_,data_stage_2__43_,
  data_stage_2__42_,data_stage_2__41_,data_stage_2__40_,data_stage_2__39_,
  data_stage_2__38_,data_stage_2__37_,data_stage_2__36_,data_stage_2__35_,data_stage_2__34_,
  data_stage_2__33_,data_stage_2__32_,data_stage_2__31_,data_stage_2__30_,
  data_stage_2__29_,data_stage_2__28_,data_stage_2__27_,data_stage_2__26_,data_stage_2__25_,
  data_stage_2__24_,data_stage_2__23_,data_stage_2__22_,data_stage_2__21_,
  data_stage_2__20_,data_stage_2__19_,data_stage_2__18_,data_stage_2__17_,data_stage_2__16_,
  data_stage_2__15_,data_stage_2__14_,data_stage_2__13_,data_stage_2__12_,
  data_stage_2__11_,data_stage_2__10_,data_stage_2__9_,data_stage_2__8_,data_stage_2__7_,
  data_stage_2__6_,data_stage_2__5_,data_stage_2__4_,data_stage_2__3_,
  data_stage_2__2_,data_stage_2__1_,data_stage_2__0_,data_stage_3__511_,data_stage_3__510_,
  data_stage_3__509_,data_stage_3__508_,data_stage_3__507_,data_stage_3__506_,
  data_stage_3__505_,data_stage_3__504_,data_stage_3__503_,data_stage_3__502_,
  data_stage_3__501_,data_stage_3__500_,data_stage_3__499_,data_stage_3__498_,
  data_stage_3__497_,data_stage_3__496_,data_stage_3__495_,data_stage_3__494_,data_stage_3__493_,
  data_stage_3__492_,data_stage_3__491_,data_stage_3__490_,data_stage_3__489_,
  data_stage_3__488_,data_stage_3__487_,data_stage_3__486_,data_stage_3__485_,
  data_stage_3__484_,data_stage_3__483_,data_stage_3__482_,data_stage_3__481_,
  data_stage_3__480_,data_stage_3__479_,data_stage_3__478_,data_stage_3__477_,data_stage_3__476_,
  data_stage_3__475_,data_stage_3__474_,data_stage_3__473_,data_stage_3__472_,
  data_stage_3__471_,data_stage_3__470_,data_stage_3__469_,data_stage_3__468_,
  data_stage_3__467_,data_stage_3__466_,data_stage_3__465_,data_stage_3__464_,
  data_stage_3__463_,data_stage_3__462_,data_stage_3__461_,data_stage_3__460_,
  data_stage_3__459_,data_stage_3__458_,data_stage_3__457_,data_stage_3__456_,data_stage_3__455_,
  data_stage_3__454_,data_stage_3__453_,data_stage_3__452_,data_stage_3__451_,
  data_stage_3__450_,data_stage_3__449_,data_stage_3__448_,data_stage_3__447_,
  data_stage_3__446_,data_stage_3__445_,data_stage_3__444_,data_stage_3__443_,
  data_stage_3__442_,data_stage_3__441_,data_stage_3__440_,data_stage_3__439_,
  data_stage_3__438_,data_stage_3__437_,data_stage_3__436_,data_stage_3__435_,data_stage_3__434_,
  data_stage_3__433_,data_stage_3__432_,data_stage_3__431_,data_stage_3__430_,
  data_stage_3__429_,data_stage_3__428_,data_stage_3__427_,data_stage_3__426_,
  data_stage_3__425_,data_stage_3__424_,data_stage_3__423_,data_stage_3__422_,
  data_stage_3__421_,data_stage_3__420_,data_stage_3__419_,data_stage_3__418_,
  data_stage_3__417_,data_stage_3__416_,data_stage_3__415_,data_stage_3__414_,data_stage_3__413_,
  data_stage_3__412_,data_stage_3__411_,data_stage_3__410_,data_stage_3__409_,
  data_stage_3__408_,data_stage_3__407_,data_stage_3__406_,data_stage_3__405_,
  data_stage_3__404_,data_stage_3__403_,data_stage_3__402_,data_stage_3__401_,
  data_stage_3__400_,data_stage_3__399_,data_stage_3__398_,data_stage_3__397_,data_stage_3__396_,
  data_stage_3__395_,data_stage_3__394_,data_stage_3__393_,data_stage_3__392_,
  data_stage_3__391_,data_stage_3__390_,data_stage_3__389_,data_stage_3__388_,
  data_stage_3__387_,data_stage_3__386_,data_stage_3__385_,data_stage_3__384_,
  data_stage_3__383_,data_stage_3__382_,data_stage_3__381_,data_stage_3__380_,
  data_stage_3__379_,data_stage_3__378_,data_stage_3__377_,data_stage_3__376_,data_stage_3__375_,
  data_stage_3__374_,data_stage_3__373_,data_stage_3__372_,data_stage_3__371_,
  data_stage_3__370_,data_stage_3__369_,data_stage_3__368_,data_stage_3__367_,
  data_stage_3__366_,data_stage_3__365_,data_stage_3__364_,data_stage_3__363_,
  data_stage_3__362_,data_stage_3__361_,data_stage_3__360_,data_stage_3__359_,
  data_stage_3__358_,data_stage_3__357_,data_stage_3__356_,data_stage_3__355_,data_stage_3__354_,
  data_stage_3__353_,data_stage_3__352_,data_stage_3__351_,data_stage_3__350_,
  data_stage_3__349_,data_stage_3__348_,data_stage_3__347_,data_stage_3__346_,
  data_stage_3__345_,data_stage_3__344_,data_stage_3__343_,data_stage_3__342_,
  data_stage_3__341_,data_stage_3__340_,data_stage_3__339_,data_stage_3__338_,
  data_stage_3__337_,data_stage_3__336_,data_stage_3__335_,data_stage_3__334_,data_stage_3__333_,
  data_stage_3__332_,data_stage_3__331_,data_stage_3__330_,data_stage_3__329_,
  data_stage_3__328_,data_stage_3__327_,data_stage_3__326_,data_stage_3__325_,
  data_stage_3__324_,data_stage_3__323_,data_stage_3__322_,data_stage_3__321_,
  data_stage_3__320_,data_stage_3__319_,data_stage_3__318_,data_stage_3__317_,data_stage_3__316_,
  data_stage_3__315_,data_stage_3__314_,data_stage_3__313_,data_stage_3__312_,
  data_stage_3__311_,data_stage_3__310_,data_stage_3__309_,data_stage_3__308_,
  data_stage_3__307_,data_stage_3__306_,data_stage_3__305_,data_stage_3__304_,
  data_stage_3__303_,data_stage_3__302_,data_stage_3__301_,data_stage_3__300_,
  data_stage_3__299_,data_stage_3__298_,data_stage_3__297_,data_stage_3__296_,data_stage_3__295_,
  data_stage_3__294_,data_stage_3__293_,data_stage_3__292_,data_stage_3__291_,
  data_stage_3__290_,data_stage_3__289_,data_stage_3__288_,data_stage_3__287_,
  data_stage_3__286_,data_stage_3__285_,data_stage_3__284_,data_stage_3__283_,
  data_stage_3__282_,data_stage_3__281_,data_stage_3__280_,data_stage_3__279_,
  data_stage_3__278_,data_stage_3__277_,data_stage_3__276_,data_stage_3__275_,data_stage_3__274_,
  data_stage_3__273_,data_stage_3__272_,data_stage_3__271_,data_stage_3__270_,
  data_stage_3__269_,data_stage_3__268_,data_stage_3__267_,data_stage_3__266_,
  data_stage_3__265_,data_stage_3__264_,data_stage_3__263_,data_stage_3__262_,
  data_stage_3__261_,data_stage_3__260_,data_stage_3__259_,data_stage_3__258_,
  data_stage_3__257_,data_stage_3__256_,data_stage_3__255_,data_stage_3__254_,data_stage_3__253_,
  data_stage_3__252_,data_stage_3__251_,data_stage_3__250_,data_stage_3__249_,
  data_stage_3__248_,data_stage_3__247_,data_stage_3__246_,data_stage_3__245_,
  data_stage_3__244_,data_stage_3__243_,data_stage_3__242_,data_stage_3__241_,
  data_stage_3__240_,data_stage_3__239_,data_stage_3__238_,data_stage_3__237_,data_stage_3__236_,
  data_stage_3__235_,data_stage_3__234_,data_stage_3__233_,data_stage_3__232_,
  data_stage_3__231_,data_stage_3__230_,data_stage_3__229_,data_stage_3__228_,
  data_stage_3__227_,data_stage_3__226_,data_stage_3__225_,data_stage_3__224_,
  data_stage_3__223_,data_stage_3__222_,data_stage_3__221_,data_stage_3__220_,
  data_stage_3__219_,data_stage_3__218_,data_stage_3__217_,data_stage_3__216_,data_stage_3__215_,
  data_stage_3__214_,data_stage_3__213_,data_stage_3__212_,data_stage_3__211_,
  data_stage_3__210_,data_stage_3__209_,data_stage_3__208_,data_stage_3__207_,
  data_stage_3__206_,data_stage_3__205_,data_stage_3__204_,data_stage_3__203_,
  data_stage_3__202_,data_stage_3__201_,data_stage_3__200_,data_stage_3__199_,
  data_stage_3__198_,data_stage_3__197_,data_stage_3__196_,data_stage_3__195_,data_stage_3__194_,
  data_stage_3__193_,data_stage_3__192_,data_stage_3__191_,data_stage_3__190_,
  data_stage_3__189_,data_stage_3__188_,data_stage_3__187_,data_stage_3__186_,
  data_stage_3__185_,data_stage_3__184_,data_stage_3__183_,data_stage_3__182_,
  data_stage_3__181_,data_stage_3__180_,data_stage_3__179_,data_stage_3__178_,
  data_stage_3__177_,data_stage_3__176_,data_stage_3__175_,data_stage_3__174_,data_stage_3__173_,
  data_stage_3__172_,data_stage_3__171_,data_stage_3__170_,data_stage_3__169_,
  data_stage_3__168_,data_stage_3__167_,data_stage_3__166_,data_stage_3__165_,
  data_stage_3__164_,data_stage_3__163_,data_stage_3__162_,data_stage_3__161_,
  data_stage_3__160_,data_stage_3__159_,data_stage_3__158_,data_stage_3__157_,data_stage_3__156_,
  data_stage_3__155_,data_stage_3__154_,data_stage_3__153_,data_stage_3__152_,
  data_stage_3__151_,data_stage_3__150_,data_stage_3__149_,data_stage_3__148_,
  data_stage_3__147_,data_stage_3__146_,data_stage_3__145_,data_stage_3__144_,
  data_stage_3__143_,data_stage_3__142_,data_stage_3__141_,data_stage_3__140_,
  data_stage_3__139_,data_stage_3__138_,data_stage_3__137_,data_stage_3__136_,data_stage_3__135_,
  data_stage_3__134_,data_stage_3__133_,data_stage_3__132_,data_stage_3__131_,
  data_stage_3__130_,data_stage_3__129_,data_stage_3__128_,data_stage_3__127_,
  data_stage_3__126_,data_stage_3__125_,data_stage_3__124_,data_stage_3__123_,
  data_stage_3__122_,data_stage_3__121_,data_stage_3__120_,data_stage_3__119_,
  data_stage_3__118_,data_stage_3__117_,data_stage_3__116_,data_stage_3__115_,data_stage_3__114_,
  data_stage_3__113_,data_stage_3__112_,data_stage_3__111_,data_stage_3__110_,
  data_stage_3__109_,data_stage_3__108_,data_stage_3__107_,data_stage_3__106_,
  data_stage_3__105_,data_stage_3__104_,data_stage_3__103_,data_stage_3__102_,
  data_stage_3__101_,data_stage_3__100_,data_stage_3__99_,data_stage_3__98_,data_stage_3__97_,
  data_stage_3__96_,data_stage_3__95_,data_stage_3__94_,data_stage_3__93_,
  data_stage_3__92_,data_stage_3__91_,data_stage_3__90_,data_stage_3__89_,data_stage_3__88_,
  data_stage_3__87_,data_stage_3__86_,data_stage_3__85_,data_stage_3__84_,
  data_stage_3__83_,data_stage_3__82_,data_stage_3__81_,data_stage_3__80_,
  data_stage_3__79_,data_stage_3__78_,data_stage_3__77_,data_stage_3__76_,data_stage_3__75_,
  data_stage_3__74_,data_stage_3__73_,data_stage_3__72_,data_stage_3__71_,
  data_stage_3__70_,data_stage_3__69_,data_stage_3__68_,data_stage_3__67_,data_stage_3__66_,
  data_stage_3__65_,data_stage_3__64_,data_stage_3__63_,data_stage_3__62_,
  data_stage_3__61_,data_stage_3__60_,data_stage_3__59_,data_stage_3__58_,data_stage_3__57_,
  data_stage_3__56_,data_stage_3__55_,data_stage_3__54_,data_stage_3__53_,
  data_stage_3__52_,data_stage_3__51_,data_stage_3__50_,data_stage_3__49_,data_stage_3__48_,
  data_stage_3__47_,data_stage_3__46_,data_stage_3__45_,data_stage_3__44_,
  data_stage_3__43_,data_stage_3__42_,data_stage_3__41_,data_stage_3__40_,
  data_stage_3__39_,data_stage_3__38_,data_stage_3__37_,data_stage_3__36_,data_stage_3__35_,
  data_stage_3__34_,data_stage_3__33_,data_stage_3__32_,data_stage_3__31_,
  data_stage_3__30_,data_stage_3__29_,data_stage_3__28_,data_stage_3__27_,data_stage_3__26_,
  data_stage_3__25_,data_stage_3__24_,data_stage_3__23_,data_stage_3__22_,
  data_stage_3__21_,data_stage_3__20_,data_stage_3__19_,data_stage_3__18_,data_stage_3__17_,
  data_stage_3__16_,data_stage_3__15_,data_stage_3__14_,data_stage_3__13_,
  data_stage_3__12_,data_stage_3__11_,data_stage_3__10_,data_stage_3__9_,data_stage_3__8_,
  data_stage_3__7_,data_stage_3__6_,data_stage_3__5_,data_stage_3__4_,
  data_stage_3__3_,data_stage_3__2_,data_stage_3__1_,data_stage_3__0_,data_stage_4__511_,
  data_stage_4__510_,data_stage_4__509_,data_stage_4__508_,data_stage_4__507_,
  data_stage_4__506_,data_stage_4__505_,data_stage_4__504_,data_stage_4__503_,
  data_stage_4__502_,data_stage_4__501_,data_stage_4__500_,data_stage_4__499_,data_stage_4__498_,
  data_stage_4__497_,data_stage_4__496_,data_stage_4__495_,data_stage_4__494_,
  data_stage_4__493_,data_stage_4__492_,data_stage_4__491_,data_stage_4__490_,
  data_stage_4__489_,data_stage_4__488_,data_stage_4__487_,data_stage_4__486_,
  data_stage_4__485_,data_stage_4__484_,data_stage_4__483_,data_stage_4__482_,
  data_stage_4__481_,data_stage_4__480_,data_stage_4__479_,data_stage_4__478_,data_stage_4__477_,
  data_stage_4__476_,data_stage_4__475_,data_stage_4__474_,data_stage_4__473_,
  data_stage_4__472_,data_stage_4__471_,data_stage_4__470_,data_stage_4__469_,
  data_stage_4__468_,data_stage_4__467_,data_stage_4__466_,data_stage_4__465_,
  data_stage_4__464_,data_stage_4__463_,data_stage_4__462_,data_stage_4__461_,
  data_stage_4__460_,data_stage_4__459_,data_stage_4__458_,data_stage_4__457_,data_stage_4__456_,
  data_stage_4__455_,data_stage_4__454_,data_stage_4__453_,data_stage_4__452_,
  data_stage_4__451_,data_stage_4__450_,data_stage_4__449_,data_stage_4__448_,
  data_stage_4__447_,data_stage_4__446_,data_stage_4__445_,data_stage_4__444_,
  data_stage_4__443_,data_stage_4__442_,data_stage_4__441_,data_stage_4__440_,
  data_stage_4__439_,data_stage_4__438_,data_stage_4__437_,data_stage_4__436_,data_stage_4__435_,
  data_stage_4__434_,data_stage_4__433_,data_stage_4__432_,data_stage_4__431_,
  data_stage_4__430_,data_stage_4__429_,data_stage_4__428_,data_stage_4__427_,
  data_stage_4__426_,data_stage_4__425_,data_stage_4__424_,data_stage_4__423_,
  data_stage_4__422_,data_stage_4__421_,data_stage_4__420_,data_stage_4__419_,data_stage_4__418_,
  data_stage_4__417_,data_stage_4__416_,data_stage_4__415_,data_stage_4__414_,
  data_stage_4__413_,data_stage_4__412_,data_stage_4__411_,data_stage_4__410_,
  data_stage_4__409_,data_stage_4__408_,data_stage_4__407_,data_stage_4__406_,
  data_stage_4__405_,data_stage_4__404_,data_stage_4__403_,data_stage_4__402_,
  data_stage_4__401_,data_stage_4__400_,data_stage_4__399_,data_stage_4__398_,data_stage_4__397_,
  data_stage_4__396_,data_stage_4__395_,data_stage_4__394_,data_stage_4__393_,
  data_stage_4__392_,data_stage_4__391_,data_stage_4__390_,data_stage_4__389_,
  data_stage_4__388_,data_stage_4__387_,data_stage_4__386_,data_stage_4__385_,
  data_stage_4__384_,data_stage_4__383_,data_stage_4__382_,data_stage_4__381_,
  data_stage_4__380_,data_stage_4__379_,data_stage_4__378_,data_stage_4__377_,data_stage_4__376_,
  data_stage_4__375_,data_stage_4__374_,data_stage_4__373_,data_stage_4__372_,
  data_stage_4__371_,data_stage_4__370_,data_stage_4__369_,data_stage_4__368_,
  data_stage_4__367_,data_stage_4__366_,data_stage_4__365_,data_stage_4__364_,
  data_stage_4__363_,data_stage_4__362_,data_stage_4__361_,data_stage_4__360_,
  data_stage_4__359_,data_stage_4__358_,data_stage_4__357_,data_stage_4__356_,data_stage_4__355_,
  data_stage_4__354_,data_stage_4__353_,data_stage_4__352_,data_stage_4__351_,
  data_stage_4__350_,data_stage_4__349_,data_stage_4__348_,data_stage_4__347_,
  data_stage_4__346_,data_stage_4__345_,data_stage_4__344_,data_stage_4__343_,
  data_stage_4__342_,data_stage_4__341_,data_stage_4__340_,data_stage_4__339_,data_stage_4__338_,
  data_stage_4__337_,data_stage_4__336_,data_stage_4__335_,data_stage_4__334_,
  data_stage_4__333_,data_stage_4__332_,data_stage_4__331_,data_stage_4__330_,
  data_stage_4__329_,data_stage_4__328_,data_stage_4__327_,data_stage_4__326_,
  data_stage_4__325_,data_stage_4__324_,data_stage_4__323_,data_stage_4__322_,
  data_stage_4__321_,data_stage_4__320_,data_stage_4__319_,data_stage_4__318_,data_stage_4__317_,
  data_stage_4__316_,data_stage_4__315_,data_stage_4__314_,data_stage_4__313_,
  data_stage_4__312_,data_stage_4__311_,data_stage_4__310_,data_stage_4__309_,
  data_stage_4__308_,data_stage_4__307_,data_stage_4__306_,data_stage_4__305_,
  data_stage_4__304_,data_stage_4__303_,data_stage_4__302_,data_stage_4__301_,
  data_stage_4__300_,data_stage_4__299_,data_stage_4__298_,data_stage_4__297_,data_stage_4__296_,
  data_stage_4__295_,data_stage_4__294_,data_stage_4__293_,data_stage_4__292_,
  data_stage_4__291_,data_stage_4__290_,data_stage_4__289_,data_stage_4__288_,
  data_stage_4__287_,data_stage_4__286_,data_stage_4__285_,data_stage_4__284_,
  data_stage_4__283_,data_stage_4__282_,data_stage_4__281_,data_stage_4__280_,
  data_stage_4__279_,data_stage_4__278_,data_stage_4__277_,data_stage_4__276_,data_stage_4__275_,
  data_stage_4__274_,data_stage_4__273_,data_stage_4__272_,data_stage_4__271_,
  data_stage_4__270_,data_stage_4__269_,data_stage_4__268_,data_stage_4__267_,
  data_stage_4__266_,data_stage_4__265_,data_stage_4__264_,data_stage_4__263_,
  data_stage_4__262_,data_stage_4__261_,data_stage_4__260_,data_stage_4__259_,data_stage_4__258_,
  data_stage_4__257_,data_stage_4__256_,data_stage_4__255_,data_stage_4__254_,
  data_stage_4__253_,data_stage_4__252_,data_stage_4__251_,data_stage_4__250_,
  data_stage_4__249_,data_stage_4__248_,data_stage_4__247_,data_stage_4__246_,
  data_stage_4__245_,data_stage_4__244_,data_stage_4__243_,data_stage_4__242_,
  data_stage_4__241_,data_stage_4__240_,data_stage_4__239_,data_stage_4__238_,data_stage_4__237_,
  data_stage_4__236_,data_stage_4__235_,data_stage_4__234_,data_stage_4__233_,
  data_stage_4__232_,data_stage_4__231_,data_stage_4__230_,data_stage_4__229_,
  data_stage_4__228_,data_stage_4__227_,data_stage_4__226_,data_stage_4__225_,
  data_stage_4__224_,data_stage_4__223_,data_stage_4__222_,data_stage_4__221_,
  data_stage_4__220_,data_stage_4__219_,data_stage_4__218_,data_stage_4__217_,data_stage_4__216_,
  data_stage_4__215_,data_stage_4__214_,data_stage_4__213_,data_stage_4__212_,
  data_stage_4__211_,data_stage_4__210_,data_stage_4__209_,data_stage_4__208_,
  data_stage_4__207_,data_stage_4__206_,data_stage_4__205_,data_stage_4__204_,
  data_stage_4__203_,data_stage_4__202_,data_stage_4__201_,data_stage_4__200_,
  data_stage_4__199_,data_stage_4__198_,data_stage_4__197_,data_stage_4__196_,data_stage_4__195_,
  data_stage_4__194_,data_stage_4__193_,data_stage_4__192_,data_stage_4__191_,
  data_stage_4__190_,data_stage_4__189_,data_stage_4__188_,data_stage_4__187_,
  data_stage_4__186_,data_stage_4__185_,data_stage_4__184_,data_stage_4__183_,
  data_stage_4__182_,data_stage_4__181_,data_stage_4__180_,data_stage_4__179_,data_stage_4__178_,
  data_stage_4__177_,data_stage_4__176_,data_stage_4__175_,data_stage_4__174_,
  data_stage_4__173_,data_stage_4__172_,data_stage_4__171_,data_stage_4__170_,
  data_stage_4__169_,data_stage_4__168_,data_stage_4__167_,data_stage_4__166_,
  data_stage_4__165_,data_stage_4__164_,data_stage_4__163_,data_stage_4__162_,
  data_stage_4__161_,data_stage_4__160_,data_stage_4__159_,data_stage_4__158_,data_stage_4__157_,
  data_stage_4__156_,data_stage_4__155_,data_stage_4__154_,data_stage_4__153_,
  data_stage_4__152_,data_stage_4__151_,data_stage_4__150_,data_stage_4__149_,
  data_stage_4__148_,data_stage_4__147_,data_stage_4__146_,data_stage_4__145_,
  data_stage_4__144_,data_stage_4__143_,data_stage_4__142_,data_stage_4__141_,
  data_stage_4__140_,data_stage_4__139_,data_stage_4__138_,data_stage_4__137_,data_stage_4__136_,
  data_stage_4__135_,data_stage_4__134_,data_stage_4__133_,data_stage_4__132_,
  data_stage_4__131_,data_stage_4__130_,data_stage_4__129_,data_stage_4__128_,
  data_stage_4__127_,data_stage_4__126_,data_stage_4__125_,data_stage_4__124_,
  data_stage_4__123_,data_stage_4__122_,data_stage_4__121_,data_stage_4__120_,
  data_stage_4__119_,data_stage_4__118_,data_stage_4__117_,data_stage_4__116_,data_stage_4__115_,
  data_stage_4__114_,data_stage_4__113_,data_stage_4__112_,data_stage_4__111_,
  data_stage_4__110_,data_stage_4__109_,data_stage_4__108_,data_stage_4__107_,
  data_stage_4__106_,data_stage_4__105_,data_stage_4__104_,data_stage_4__103_,
  data_stage_4__102_,data_stage_4__101_,data_stage_4__100_,data_stage_4__99_,data_stage_4__98_,
  data_stage_4__97_,data_stage_4__96_,data_stage_4__95_,data_stage_4__94_,
  data_stage_4__93_,data_stage_4__92_,data_stage_4__91_,data_stage_4__90_,data_stage_4__89_,
  data_stage_4__88_,data_stage_4__87_,data_stage_4__86_,data_stage_4__85_,
  data_stage_4__84_,data_stage_4__83_,data_stage_4__82_,data_stage_4__81_,
  data_stage_4__80_,data_stage_4__79_,data_stage_4__78_,data_stage_4__77_,data_stage_4__76_,
  data_stage_4__75_,data_stage_4__74_,data_stage_4__73_,data_stage_4__72_,
  data_stage_4__71_,data_stage_4__70_,data_stage_4__69_,data_stage_4__68_,data_stage_4__67_,
  data_stage_4__66_,data_stage_4__65_,data_stage_4__64_,data_stage_4__63_,
  data_stage_4__62_,data_stage_4__61_,data_stage_4__60_,data_stage_4__59_,data_stage_4__58_,
  data_stage_4__57_,data_stage_4__56_,data_stage_4__55_,data_stage_4__54_,
  data_stage_4__53_,data_stage_4__52_,data_stage_4__51_,data_stage_4__50_,data_stage_4__49_,
  data_stage_4__48_,data_stage_4__47_,data_stage_4__46_,data_stage_4__45_,
  data_stage_4__44_,data_stage_4__43_,data_stage_4__42_,data_stage_4__41_,
  data_stage_4__40_,data_stage_4__39_,data_stage_4__38_,data_stage_4__37_,data_stage_4__36_,
  data_stage_4__35_,data_stage_4__34_,data_stage_4__33_,data_stage_4__32_,
  data_stage_4__31_,data_stage_4__30_,data_stage_4__29_,data_stage_4__28_,data_stage_4__27_,
  data_stage_4__26_,data_stage_4__25_,data_stage_4__24_,data_stage_4__23_,
  data_stage_4__22_,data_stage_4__21_,data_stage_4__20_,data_stage_4__19_,data_stage_4__18_,
  data_stage_4__17_,data_stage_4__16_,data_stage_4__15_,data_stage_4__14_,
  data_stage_4__13_,data_stage_4__12_,data_stage_4__11_,data_stage_4__10_,data_stage_4__9_,
  data_stage_4__8_,data_stage_4__7_,data_stage_4__6_,data_stage_4__5_,
  data_stage_4__4_,data_stage_4__3_,data_stage_4__2_,data_stage_4__1_,data_stage_4__0_;

  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_0_.swap_inst 
  (
    .data_i(data_i[31:0]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_1_.swap_inst 
  (
    .data_i(data_i[63:32]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_2_.swap_inst 
  (
    .data_i(data_i[95:64]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_3_.swap_inst 
  (
    .data_i(data_i[127:96]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_4_.swap_inst 
  (
    .data_i(data_i[159:128]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_5_.swap_inst 
  (
    .data_i(data_i[191:160]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_6_.swap_inst 
  (
    .data_i(data_i[223:192]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_7_.swap_inst 
  (
    .data_i(data_i[255:224]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_8_.swap_inst 
  (
    .data_i(data_i[287:256]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_9_.swap_inst 
  (
    .data_i(data_i[319:288]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_10_.swap_inst 
  (
    .data_i(data_i[351:320]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_11_.swap_inst 
  (
    .data_i(data_i[383:352]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_12_.swap_inst 
  (
    .data_i(data_i[415:384]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_13_.swap_inst 
  (
    .data_i(data_i[447:416]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_14_.swap_inst 
  (
    .data_i(data_i[479:448]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_ })
  );


  bsg_swap_width_p16
  \mux_stage_0_.mux_swap_15_.swap_inst 
  (
    .data_i(data_i[511:480]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_ })
  );


  bsg_swap_width_p32
  \mux_stage_1_.mux_swap_0_.swap_inst 
  (
    .data_i({ data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ })
  );


  bsg_swap_width_p32
  \mux_stage_1_.mux_swap_1_.swap_inst 
  (
    .data_i({ data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_ })
  );


  bsg_swap_width_p32
  \mux_stage_1_.mux_swap_2_.swap_inst 
  (
    .data_i({ data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_ })
  );


  bsg_swap_width_p32
  \mux_stage_1_.mux_swap_3_.swap_inst 
  (
    .data_i({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_ })
  );


  bsg_swap_width_p32
  \mux_stage_1_.mux_swap_4_.swap_inst 
  (
    .data_i({ data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_ })
  );


  bsg_swap_width_p32
  \mux_stage_1_.mux_swap_5_.swap_inst 
  (
    .data_i({ data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_ })
  );


  bsg_swap_width_p32
  \mux_stage_1_.mux_swap_6_.swap_inst 
  (
    .data_i({ data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_ })
  );


  bsg_swap_width_p32
  \mux_stage_1_.mux_swap_7_.swap_inst 
  (
    .data_i({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_ })
  );


  bsg_swap_width_p64
  \mux_stage_2_.mux_swap_0_.swap_inst 
  (
    .data_i({ data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__127_, data_stage_3__126_, data_stage_3__125_, data_stage_3__124_, data_stage_3__123_, data_stage_3__122_, data_stage_3__121_, data_stage_3__120_, data_stage_3__119_, data_stage_3__118_, data_stage_3__117_, data_stage_3__116_, data_stage_3__115_, data_stage_3__114_, data_stage_3__113_, data_stage_3__112_, data_stage_3__111_, data_stage_3__110_, data_stage_3__109_, data_stage_3__108_, data_stage_3__107_, data_stage_3__106_, data_stage_3__105_, data_stage_3__104_, data_stage_3__103_, data_stage_3__102_, data_stage_3__101_, data_stage_3__100_, data_stage_3__99_, data_stage_3__98_, data_stage_3__97_, data_stage_3__96_, data_stage_3__95_, data_stage_3__94_, data_stage_3__93_, data_stage_3__92_, data_stage_3__91_, data_stage_3__90_, data_stage_3__89_, data_stage_3__88_, data_stage_3__87_, data_stage_3__86_, data_stage_3__85_, data_stage_3__84_, data_stage_3__83_, data_stage_3__82_, data_stage_3__81_, data_stage_3__80_, data_stage_3__79_, data_stage_3__78_, data_stage_3__77_, data_stage_3__76_, data_stage_3__75_, data_stage_3__74_, data_stage_3__73_, data_stage_3__72_, data_stage_3__71_, data_stage_3__70_, data_stage_3__69_, data_stage_3__68_, data_stage_3__67_, data_stage_3__66_, data_stage_3__65_, data_stage_3__64_, data_stage_3__63_, data_stage_3__62_, data_stage_3__61_, data_stage_3__60_, data_stage_3__59_, data_stage_3__58_, data_stage_3__57_, data_stage_3__56_, data_stage_3__55_, data_stage_3__54_, data_stage_3__53_, data_stage_3__52_, data_stage_3__51_, data_stage_3__50_, data_stage_3__49_, data_stage_3__48_, data_stage_3__47_, data_stage_3__46_, data_stage_3__45_, data_stage_3__44_, data_stage_3__43_, data_stage_3__42_, data_stage_3__41_, data_stage_3__40_, data_stage_3__39_, data_stage_3__38_, data_stage_3__37_, data_stage_3__36_, data_stage_3__35_, data_stage_3__34_, data_stage_3__33_, data_stage_3__32_, data_stage_3__31_, data_stage_3__30_, data_stage_3__29_, data_stage_3__28_, data_stage_3__27_, data_stage_3__26_, data_stage_3__25_, data_stage_3__24_, data_stage_3__23_, data_stage_3__22_, data_stage_3__21_, data_stage_3__20_, data_stage_3__19_, data_stage_3__18_, data_stage_3__17_, data_stage_3__16_, data_stage_3__15_, data_stage_3__14_, data_stage_3__13_, data_stage_3__12_, data_stage_3__11_, data_stage_3__10_, data_stage_3__9_, data_stage_3__8_, data_stage_3__7_, data_stage_3__6_, data_stage_3__5_, data_stage_3__4_, data_stage_3__3_, data_stage_3__2_, data_stage_3__1_, data_stage_3__0_ })
  );


  bsg_swap_width_p64
  \mux_stage_2_.mux_swap_1_.swap_inst 
  (
    .data_i({ data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__255_, data_stage_3__254_, data_stage_3__253_, data_stage_3__252_, data_stage_3__251_, data_stage_3__250_, data_stage_3__249_, data_stage_3__248_, data_stage_3__247_, data_stage_3__246_, data_stage_3__245_, data_stage_3__244_, data_stage_3__243_, data_stage_3__242_, data_stage_3__241_, data_stage_3__240_, data_stage_3__239_, data_stage_3__238_, data_stage_3__237_, data_stage_3__236_, data_stage_3__235_, data_stage_3__234_, data_stage_3__233_, data_stage_3__232_, data_stage_3__231_, data_stage_3__230_, data_stage_3__229_, data_stage_3__228_, data_stage_3__227_, data_stage_3__226_, data_stage_3__225_, data_stage_3__224_, data_stage_3__223_, data_stage_3__222_, data_stage_3__221_, data_stage_3__220_, data_stage_3__219_, data_stage_3__218_, data_stage_3__217_, data_stage_3__216_, data_stage_3__215_, data_stage_3__214_, data_stage_3__213_, data_stage_3__212_, data_stage_3__211_, data_stage_3__210_, data_stage_3__209_, data_stage_3__208_, data_stage_3__207_, data_stage_3__206_, data_stage_3__205_, data_stage_3__204_, data_stage_3__203_, data_stage_3__202_, data_stage_3__201_, data_stage_3__200_, data_stage_3__199_, data_stage_3__198_, data_stage_3__197_, data_stage_3__196_, data_stage_3__195_, data_stage_3__194_, data_stage_3__193_, data_stage_3__192_, data_stage_3__191_, data_stage_3__190_, data_stage_3__189_, data_stage_3__188_, data_stage_3__187_, data_stage_3__186_, data_stage_3__185_, data_stage_3__184_, data_stage_3__183_, data_stage_3__182_, data_stage_3__181_, data_stage_3__180_, data_stage_3__179_, data_stage_3__178_, data_stage_3__177_, data_stage_3__176_, data_stage_3__175_, data_stage_3__174_, data_stage_3__173_, data_stage_3__172_, data_stage_3__171_, data_stage_3__170_, data_stage_3__169_, data_stage_3__168_, data_stage_3__167_, data_stage_3__166_, data_stage_3__165_, data_stage_3__164_, data_stage_3__163_, data_stage_3__162_, data_stage_3__161_, data_stage_3__160_, data_stage_3__159_, data_stage_3__158_, data_stage_3__157_, data_stage_3__156_, data_stage_3__155_, data_stage_3__154_, data_stage_3__153_, data_stage_3__152_, data_stage_3__151_, data_stage_3__150_, data_stage_3__149_, data_stage_3__148_, data_stage_3__147_, data_stage_3__146_, data_stage_3__145_, data_stage_3__144_, data_stage_3__143_, data_stage_3__142_, data_stage_3__141_, data_stage_3__140_, data_stage_3__139_, data_stage_3__138_, data_stage_3__137_, data_stage_3__136_, data_stage_3__135_, data_stage_3__134_, data_stage_3__133_, data_stage_3__132_, data_stage_3__131_, data_stage_3__130_, data_stage_3__129_, data_stage_3__128_ })
  );


  bsg_swap_width_p64
  \mux_stage_2_.mux_swap_2_.swap_inst 
  (
    .data_i({ data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__383_, data_stage_3__382_, data_stage_3__381_, data_stage_3__380_, data_stage_3__379_, data_stage_3__378_, data_stage_3__377_, data_stage_3__376_, data_stage_3__375_, data_stage_3__374_, data_stage_3__373_, data_stage_3__372_, data_stage_3__371_, data_stage_3__370_, data_stage_3__369_, data_stage_3__368_, data_stage_3__367_, data_stage_3__366_, data_stage_3__365_, data_stage_3__364_, data_stage_3__363_, data_stage_3__362_, data_stage_3__361_, data_stage_3__360_, data_stage_3__359_, data_stage_3__358_, data_stage_3__357_, data_stage_3__356_, data_stage_3__355_, data_stage_3__354_, data_stage_3__353_, data_stage_3__352_, data_stage_3__351_, data_stage_3__350_, data_stage_3__349_, data_stage_3__348_, data_stage_3__347_, data_stage_3__346_, data_stage_3__345_, data_stage_3__344_, data_stage_3__343_, data_stage_3__342_, data_stage_3__341_, data_stage_3__340_, data_stage_3__339_, data_stage_3__338_, data_stage_3__337_, data_stage_3__336_, data_stage_3__335_, data_stage_3__334_, data_stage_3__333_, data_stage_3__332_, data_stage_3__331_, data_stage_3__330_, data_stage_3__329_, data_stage_3__328_, data_stage_3__327_, data_stage_3__326_, data_stage_3__325_, data_stage_3__324_, data_stage_3__323_, data_stage_3__322_, data_stage_3__321_, data_stage_3__320_, data_stage_3__319_, data_stage_3__318_, data_stage_3__317_, data_stage_3__316_, data_stage_3__315_, data_stage_3__314_, data_stage_3__313_, data_stage_3__312_, data_stage_3__311_, data_stage_3__310_, data_stage_3__309_, data_stage_3__308_, data_stage_3__307_, data_stage_3__306_, data_stage_3__305_, data_stage_3__304_, data_stage_3__303_, data_stage_3__302_, data_stage_3__301_, data_stage_3__300_, data_stage_3__299_, data_stage_3__298_, data_stage_3__297_, data_stage_3__296_, data_stage_3__295_, data_stage_3__294_, data_stage_3__293_, data_stage_3__292_, data_stage_3__291_, data_stage_3__290_, data_stage_3__289_, data_stage_3__288_, data_stage_3__287_, data_stage_3__286_, data_stage_3__285_, data_stage_3__284_, data_stage_3__283_, data_stage_3__282_, data_stage_3__281_, data_stage_3__280_, data_stage_3__279_, data_stage_3__278_, data_stage_3__277_, data_stage_3__276_, data_stage_3__275_, data_stage_3__274_, data_stage_3__273_, data_stage_3__272_, data_stage_3__271_, data_stage_3__270_, data_stage_3__269_, data_stage_3__268_, data_stage_3__267_, data_stage_3__266_, data_stage_3__265_, data_stage_3__264_, data_stage_3__263_, data_stage_3__262_, data_stage_3__261_, data_stage_3__260_, data_stage_3__259_, data_stage_3__258_, data_stage_3__257_, data_stage_3__256_ })
  );


  bsg_swap_width_p64
  \mux_stage_2_.mux_swap_3_.swap_inst 
  (
    .data_i({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__511_, data_stage_3__510_, data_stage_3__509_, data_stage_3__508_, data_stage_3__507_, data_stage_3__506_, data_stage_3__505_, data_stage_3__504_, data_stage_3__503_, data_stage_3__502_, data_stage_3__501_, data_stage_3__500_, data_stage_3__499_, data_stage_3__498_, data_stage_3__497_, data_stage_3__496_, data_stage_3__495_, data_stage_3__494_, data_stage_3__493_, data_stage_3__492_, data_stage_3__491_, data_stage_3__490_, data_stage_3__489_, data_stage_3__488_, data_stage_3__487_, data_stage_3__486_, data_stage_3__485_, data_stage_3__484_, data_stage_3__483_, data_stage_3__482_, data_stage_3__481_, data_stage_3__480_, data_stage_3__479_, data_stage_3__478_, data_stage_3__477_, data_stage_3__476_, data_stage_3__475_, data_stage_3__474_, data_stage_3__473_, data_stage_3__472_, data_stage_3__471_, data_stage_3__470_, data_stage_3__469_, data_stage_3__468_, data_stage_3__467_, data_stage_3__466_, data_stage_3__465_, data_stage_3__464_, data_stage_3__463_, data_stage_3__462_, data_stage_3__461_, data_stage_3__460_, data_stage_3__459_, data_stage_3__458_, data_stage_3__457_, data_stage_3__456_, data_stage_3__455_, data_stage_3__454_, data_stage_3__453_, data_stage_3__452_, data_stage_3__451_, data_stage_3__450_, data_stage_3__449_, data_stage_3__448_, data_stage_3__447_, data_stage_3__446_, data_stage_3__445_, data_stage_3__444_, data_stage_3__443_, data_stage_3__442_, data_stage_3__441_, data_stage_3__440_, data_stage_3__439_, data_stage_3__438_, data_stage_3__437_, data_stage_3__436_, data_stage_3__435_, data_stage_3__434_, data_stage_3__433_, data_stage_3__432_, data_stage_3__431_, data_stage_3__430_, data_stage_3__429_, data_stage_3__428_, data_stage_3__427_, data_stage_3__426_, data_stage_3__425_, data_stage_3__424_, data_stage_3__423_, data_stage_3__422_, data_stage_3__421_, data_stage_3__420_, data_stage_3__419_, data_stage_3__418_, data_stage_3__417_, data_stage_3__416_, data_stage_3__415_, data_stage_3__414_, data_stage_3__413_, data_stage_3__412_, data_stage_3__411_, data_stage_3__410_, data_stage_3__409_, data_stage_3__408_, data_stage_3__407_, data_stage_3__406_, data_stage_3__405_, data_stage_3__404_, data_stage_3__403_, data_stage_3__402_, data_stage_3__401_, data_stage_3__400_, data_stage_3__399_, data_stage_3__398_, data_stage_3__397_, data_stage_3__396_, data_stage_3__395_, data_stage_3__394_, data_stage_3__393_, data_stage_3__392_, data_stage_3__391_, data_stage_3__390_, data_stage_3__389_, data_stage_3__388_, data_stage_3__387_, data_stage_3__386_, data_stage_3__385_, data_stage_3__384_ })
  );


  bsg_swap_width_p128
  \mux_stage_3_.mux_swap_0_.swap_inst 
  (
    .data_i({ data_stage_3__255_, data_stage_3__254_, data_stage_3__253_, data_stage_3__252_, data_stage_3__251_, data_stage_3__250_, data_stage_3__249_, data_stage_3__248_, data_stage_3__247_, data_stage_3__246_, data_stage_3__245_, data_stage_3__244_, data_stage_3__243_, data_stage_3__242_, data_stage_3__241_, data_stage_3__240_, data_stage_3__239_, data_stage_3__238_, data_stage_3__237_, data_stage_3__236_, data_stage_3__235_, data_stage_3__234_, data_stage_3__233_, data_stage_3__232_, data_stage_3__231_, data_stage_3__230_, data_stage_3__229_, data_stage_3__228_, data_stage_3__227_, data_stage_3__226_, data_stage_3__225_, data_stage_3__224_, data_stage_3__223_, data_stage_3__222_, data_stage_3__221_, data_stage_3__220_, data_stage_3__219_, data_stage_3__218_, data_stage_3__217_, data_stage_3__216_, data_stage_3__215_, data_stage_3__214_, data_stage_3__213_, data_stage_3__212_, data_stage_3__211_, data_stage_3__210_, data_stage_3__209_, data_stage_3__208_, data_stage_3__207_, data_stage_3__206_, data_stage_3__205_, data_stage_3__204_, data_stage_3__203_, data_stage_3__202_, data_stage_3__201_, data_stage_3__200_, data_stage_3__199_, data_stage_3__198_, data_stage_3__197_, data_stage_3__196_, data_stage_3__195_, data_stage_3__194_, data_stage_3__193_, data_stage_3__192_, data_stage_3__191_, data_stage_3__190_, data_stage_3__189_, data_stage_3__188_, data_stage_3__187_, data_stage_3__186_, data_stage_3__185_, data_stage_3__184_, data_stage_3__183_, data_stage_3__182_, data_stage_3__181_, data_stage_3__180_, data_stage_3__179_, data_stage_3__178_, data_stage_3__177_, data_stage_3__176_, data_stage_3__175_, data_stage_3__174_, data_stage_3__173_, data_stage_3__172_, data_stage_3__171_, data_stage_3__170_, data_stage_3__169_, data_stage_3__168_, data_stage_3__167_, data_stage_3__166_, data_stage_3__165_, data_stage_3__164_, data_stage_3__163_, data_stage_3__162_, data_stage_3__161_, data_stage_3__160_, data_stage_3__159_, data_stage_3__158_, data_stage_3__157_, data_stage_3__156_, data_stage_3__155_, data_stage_3__154_, data_stage_3__153_, data_stage_3__152_, data_stage_3__151_, data_stage_3__150_, data_stage_3__149_, data_stage_3__148_, data_stage_3__147_, data_stage_3__146_, data_stage_3__145_, data_stage_3__144_, data_stage_3__143_, data_stage_3__142_, data_stage_3__141_, data_stage_3__140_, data_stage_3__139_, data_stage_3__138_, data_stage_3__137_, data_stage_3__136_, data_stage_3__135_, data_stage_3__134_, data_stage_3__133_, data_stage_3__132_, data_stage_3__131_, data_stage_3__130_, data_stage_3__129_, data_stage_3__128_, data_stage_3__127_, data_stage_3__126_, data_stage_3__125_, data_stage_3__124_, data_stage_3__123_, data_stage_3__122_, data_stage_3__121_, data_stage_3__120_, data_stage_3__119_, data_stage_3__118_, data_stage_3__117_, data_stage_3__116_, data_stage_3__115_, data_stage_3__114_, data_stage_3__113_, data_stage_3__112_, data_stage_3__111_, data_stage_3__110_, data_stage_3__109_, data_stage_3__108_, data_stage_3__107_, data_stage_3__106_, data_stage_3__105_, data_stage_3__104_, data_stage_3__103_, data_stage_3__102_, data_stage_3__101_, data_stage_3__100_, data_stage_3__99_, data_stage_3__98_, data_stage_3__97_, data_stage_3__96_, data_stage_3__95_, data_stage_3__94_, data_stage_3__93_, data_stage_3__92_, data_stage_3__91_, data_stage_3__90_, data_stage_3__89_, data_stage_3__88_, data_stage_3__87_, data_stage_3__86_, data_stage_3__85_, data_stage_3__84_, data_stage_3__83_, data_stage_3__82_, data_stage_3__81_, data_stage_3__80_, data_stage_3__79_, data_stage_3__78_, data_stage_3__77_, data_stage_3__76_, data_stage_3__75_, data_stage_3__74_, data_stage_3__73_, data_stage_3__72_, data_stage_3__71_, data_stage_3__70_, data_stage_3__69_, data_stage_3__68_, data_stage_3__67_, data_stage_3__66_, data_stage_3__65_, data_stage_3__64_, data_stage_3__63_, data_stage_3__62_, data_stage_3__61_, data_stage_3__60_, data_stage_3__59_, data_stage_3__58_, data_stage_3__57_, data_stage_3__56_, data_stage_3__55_, data_stage_3__54_, data_stage_3__53_, data_stage_3__52_, data_stage_3__51_, data_stage_3__50_, data_stage_3__49_, data_stage_3__48_, data_stage_3__47_, data_stage_3__46_, data_stage_3__45_, data_stage_3__44_, data_stage_3__43_, data_stage_3__42_, data_stage_3__41_, data_stage_3__40_, data_stage_3__39_, data_stage_3__38_, data_stage_3__37_, data_stage_3__36_, data_stage_3__35_, data_stage_3__34_, data_stage_3__33_, data_stage_3__32_, data_stage_3__31_, data_stage_3__30_, data_stage_3__29_, data_stage_3__28_, data_stage_3__27_, data_stage_3__26_, data_stage_3__25_, data_stage_3__24_, data_stage_3__23_, data_stage_3__22_, data_stage_3__21_, data_stage_3__20_, data_stage_3__19_, data_stage_3__18_, data_stage_3__17_, data_stage_3__16_, data_stage_3__15_, data_stage_3__14_, data_stage_3__13_, data_stage_3__12_, data_stage_3__11_, data_stage_3__10_, data_stage_3__9_, data_stage_3__8_, data_stage_3__7_, data_stage_3__6_, data_stage_3__5_, data_stage_3__4_, data_stage_3__3_, data_stage_3__2_, data_stage_3__1_, data_stage_3__0_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__255_, data_stage_4__254_, data_stage_4__253_, data_stage_4__252_, data_stage_4__251_, data_stage_4__250_, data_stage_4__249_, data_stage_4__248_, data_stage_4__247_, data_stage_4__246_, data_stage_4__245_, data_stage_4__244_, data_stage_4__243_, data_stage_4__242_, data_stage_4__241_, data_stage_4__240_, data_stage_4__239_, data_stage_4__238_, data_stage_4__237_, data_stage_4__236_, data_stage_4__235_, data_stage_4__234_, data_stage_4__233_, data_stage_4__232_, data_stage_4__231_, data_stage_4__230_, data_stage_4__229_, data_stage_4__228_, data_stage_4__227_, data_stage_4__226_, data_stage_4__225_, data_stage_4__224_, data_stage_4__223_, data_stage_4__222_, data_stage_4__221_, data_stage_4__220_, data_stage_4__219_, data_stage_4__218_, data_stage_4__217_, data_stage_4__216_, data_stage_4__215_, data_stage_4__214_, data_stage_4__213_, data_stage_4__212_, data_stage_4__211_, data_stage_4__210_, data_stage_4__209_, data_stage_4__208_, data_stage_4__207_, data_stage_4__206_, data_stage_4__205_, data_stage_4__204_, data_stage_4__203_, data_stage_4__202_, data_stage_4__201_, data_stage_4__200_, data_stage_4__199_, data_stage_4__198_, data_stage_4__197_, data_stage_4__196_, data_stage_4__195_, data_stage_4__194_, data_stage_4__193_, data_stage_4__192_, data_stage_4__191_, data_stage_4__190_, data_stage_4__189_, data_stage_4__188_, data_stage_4__187_, data_stage_4__186_, data_stage_4__185_, data_stage_4__184_, data_stage_4__183_, data_stage_4__182_, data_stage_4__181_, data_stage_4__180_, data_stage_4__179_, data_stage_4__178_, data_stage_4__177_, data_stage_4__176_, data_stage_4__175_, data_stage_4__174_, data_stage_4__173_, data_stage_4__172_, data_stage_4__171_, data_stage_4__170_, data_stage_4__169_, data_stage_4__168_, data_stage_4__167_, data_stage_4__166_, data_stage_4__165_, data_stage_4__164_, data_stage_4__163_, data_stage_4__162_, data_stage_4__161_, data_stage_4__160_, data_stage_4__159_, data_stage_4__158_, data_stage_4__157_, data_stage_4__156_, data_stage_4__155_, data_stage_4__154_, data_stage_4__153_, data_stage_4__152_, data_stage_4__151_, data_stage_4__150_, data_stage_4__149_, data_stage_4__148_, data_stage_4__147_, data_stage_4__146_, data_stage_4__145_, data_stage_4__144_, data_stage_4__143_, data_stage_4__142_, data_stage_4__141_, data_stage_4__140_, data_stage_4__139_, data_stage_4__138_, data_stage_4__137_, data_stage_4__136_, data_stage_4__135_, data_stage_4__134_, data_stage_4__133_, data_stage_4__132_, data_stage_4__131_, data_stage_4__130_, data_stage_4__129_, data_stage_4__128_, data_stage_4__127_, data_stage_4__126_, data_stage_4__125_, data_stage_4__124_, data_stage_4__123_, data_stage_4__122_, data_stage_4__121_, data_stage_4__120_, data_stage_4__119_, data_stage_4__118_, data_stage_4__117_, data_stage_4__116_, data_stage_4__115_, data_stage_4__114_, data_stage_4__113_, data_stage_4__112_, data_stage_4__111_, data_stage_4__110_, data_stage_4__109_, data_stage_4__108_, data_stage_4__107_, data_stage_4__106_, data_stage_4__105_, data_stage_4__104_, data_stage_4__103_, data_stage_4__102_, data_stage_4__101_, data_stage_4__100_, data_stage_4__99_, data_stage_4__98_, data_stage_4__97_, data_stage_4__96_, data_stage_4__95_, data_stage_4__94_, data_stage_4__93_, data_stage_4__92_, data_stage_4__91_, data_stage_4__90_, data_stage_4__89_, data_stage_4__88_, data_stage_4__87_, data_stage_4__86_, data_stage_4__85_, data_stage_4__84_, data_stage_4__83_, data_stage_4__82_, data_stage_4__81_, data_stage_4__80_, data_stage_4__79_, data_stage_4__78_, data_stage_4__77_, data_stage_4__76_, data_stage_4__75_, data_stage_4__74_, data_stage_4__73_, data_stage_4__72_, data_stage_4__71_, data_stage_4__70_, data_stage_4__69_, data_stage_4__68_, data_stage_4__67_, data_stage_4__66_, data_stage_4__65_, data_stage_4__64_, data_stage_4__63_, data_stage_4__62_, data_stage_4__61_, data_stage_4__60_, data_stage_4__59_, data_stage_4__58_, data_stage_4__57_, data_stage_4__56_, data_stage_4__55_, data_stage_4__54_, data_stage_4__53_, data_stage_4__52_, data_stage_4__51_, data_stage_4__50_, data_stage_4__49_, data_stage_4__48_, data_stage_4__47_, data_stage_4__46_, data_stage_4__45_, data_stage_4__44_, data_stage_4__43_, data_stage_4__42_, data_stage_4__41_, data_stage_4__40_, data_stage_4__39_, data_stage_4__38_, data_stage_4__37_, data_stage_4__36_, data_stage_4__35_, data_stage_4__34_, data_stage_4__33_, data_stage_4__32_, data_stage_4__31_, data_stage_4__30_, data_stage_4__29_, data_stage_4__28_, data_stage_4__27_, data_stage_4__26_, data_stage_4__25_, data_stage_4__24_, data_stage_4__23_, data_stage_4__22_, data_stage_4__21_, data_stage_4__20_, data_stage_4__19_, data_stage_4__18_, data_stage_4__17_, data_stage_4__16_, data_stage_4__15_, data_stage_4__14_, data_stage_4__13_, data_stage_4__12_, data_stage_4__11_, data_stage_4__10_, data_stage_4__9_, data_stage_4__8_, data_stage_4__7_, data_stage_4__6_, data_stage_4__5_, data_stage_4__4_, data_stage_4__3_, data_stage_4__2_, data_stage_4__1_, data_stage_4__0_ })
  );


  bsg_swap_width_p128
  \mux_stage_3_.mux_swap_1_.swap_inst 
  (
    .data_i({ data_stage_3__511_, data_stage_3__510_, data_stage_3__509_, data_stage_3__508_, data_stage_3__507_, data_stage_3__506_, data_stage_3__505_, data_stage_3__504_, data_stage_3__503_, data_stage_3__502_, data_stage_3__501_, data_stage_3__500_, data_stage_3__499_, data_stage_3__498_, data_stage_3__497_, data_stage_3__496_, data_stage_3__495_, data_stage_3__494_, data_stage_3__493_, data_stage_3__492_, data_stage_3__491_, data_stage_3__490_, data_stage_3__489_, data_stage_3__488_, data_stage_3__487_, data_stage_3__486_, data_stage_3__485_, data_stage_3__484_, data_stage_3__483_, data_stage_3__482_, data_stage_3__481_, data_stage_3__480_, data_stage_3__479_, data_stage_3__478_, data_stage_3__477_, data_stage_3__476_, data_stage_3__475_, data_stage_3__474_, data_stage_3__473_, data_stage_3__472_, data_stage_3__471_, data_stage_3__470_, data_stage_3__469_, data_stage_3__468_, data_stage_3__467_, data_stage_3__466_, data_stage_3__465_, data_stage_3__464_, data_stage_3__463_, data_stage_3__462_, data_stage_3__461_, data_stage_3__460_, data_stage_3__459_, data_stage_3__458_, data_stage_3__457_, data_stage_3__456_, data_stage_3__455_, data_stage_3__454_, data_stage_3__453_, data_stage_3__452_, data_stage_3__451_, data_stage_3__450_, data_stage_3__449_, data_stage_3__448_, data_stage_3__447_, data_stage_3__446_, data_stage_3__445_, data_stage_3__444_, data_stage_3__443_, data_stage_3__442_, data_stage_3__441_, data_stage_3__440_, data_stage_3__439_, data_stage_3__438_, data_stage_3__437_, data_stage_3__436_, data_stage_3__435_, data_stage_3__434_, data_stage_3__433_, data_stage_3__432_, data_stage_3__431_, data_stage_3__430_, data_stage_3__429_, data_stage_3__428_, data_stage_3__427_, data_stage_3__426_, data_stage_3__425_, data_stage_3__424_, data_stage_3__423_, data_stage_3__422_, data_stage_3__421_, data_stage_3__420_, data_stage_3__419_, data_stage_3__418_, data_stage_3__417_, data_stage_3__416_, data_stage_3__415_, data_stage_3__414_, data_stage_3__413_, data_stage_3__412_, data_stage_3__411_, data_stage_3__410_, data_stage_3__409_, data_stage_3__408_, data_stage_3__407_, data_stage_3__406_, data_stage_3__405_, data_stage_3__404_, data_stage_3__403_, data_stage_3__402_, data_stage_3__401_, data_stage_3__400_, data_stage_3__399_, data_stage_3__398_, data_stage_3__397_, data_stage_3__396_, data_stage_3__395_, data_stage_3__394_, data_stage_3__393_, data_stage_3__392_, data_stage_3__391_, data_stage_3__390_, data_stage_3__389_, data_stage_3__388_, data_stage_3__387_, data_stage_3__386_, data_stage_3__385_, data_stage_3__384_, data_stage_3__383_, data_stage_3__382_, data_stage_3__381_, data_stage_3__380_, data_stage_3__379_, data_stage_3__378_, data_stage_3__377_, data_stage_3__376_, data_stage_3__375_, data_stage_3__374_, data_stage_3__373_, data_stage_3__372_, data_stage_3__371_, data_stage_3__370_, data_stage_3__369_, data_stage_3__368_, data_stage_3__367_, data_stage_3__366_, data_stage_3__365_, data_stage_3__364_, data_stage_3__363_, data_stage_3__362_, data_stage_3__361_, data_stage_3__360_, data_stage_3__359_, data_stage_3__358_, data_stage_3__357_, data_stage_3__356_, data_stage_3__355_, data_stage_3__354_, data_stage_3__353_, data_stage_3__352_, data_stage_3__351_, data_stage_3__350_, data_stage_3__349_, data_stage_3__348_, data_stage_3__347_, data_stage_3__346_, data_stage_3__345_, data_stage_3__344_, data_stage_3__343_, data_stage_3__342_, data_stage_3__341_, data_stage_3__340_, data_stage_3__339_, data_stage_3__338_, data_stage_3__337_, data_stage_3__336_, data_stage_3__335_, data_stage_3__334_, data_stage_3__333_, data_stage_3__332_, data_stage_3__331_, data_stage_3__330_, data_stage_3__329_, data_stage_3__328_, data_stage_3__327_, data_stage_3__326_, data_stage_3__325_, data_stage_3__324_, data_stage_3__323_, data_stage_3__322_, data_stage_3__321_, data_stage_3__320_, data_stage_3__319_, data_stage_3__318_, data_stage_3__317_, data_stage_3__316_, data_stage_3__315_, data_stage_3__314_, data_stage_3__313_, data_stage_3__312_, data_stage_3__311_, data_stage_3__310_, data_stage_3__309_, data_stage_3__308_, data_stage_3__307_, data_stage_3__306_, data_stage_3__305_, data_stage_3__304_, data_stage_3__303_, data_stage_3__302_, data_stage_3__301_, data_stage_3__300_, data_stage_3__299_, data_stage_3__298_, data_stage_3__297_, data_stage_3__296_, data_stage_3__295_, data_stage_3__294_, data_stage_3__293_, data_stage_3__292_, data_stage_3__291_, data_stage_3__290_, data_stage_3__289_, data_stage_3__288_, data_stage_3__287_, data_stage_3__286_, data_stage_3__285_, data_stage_3__284_, data_stage_3__283_, data_stage_3__282_, data_stage_3__281_, data_stage_3__280_, data_stage_3__279_, data_stage_3__278_, data_stage_3__277_, data_stage_3__276_, data_stage_3__275_, data_stage_3__274_, data_stage_3__273_, data_stage_3__272_, data_stage_3__271_, data_stage_3__270_, data_stage_3__269_, data_stage_3__268_, data_stage_3__267_, data_stage_3__266_, data_stage_3__265_, data_stage_3__264_, data_stage_3__263_, data_stage_3__262_, data_stage_3__261_, data_stage_3__260_, data_stage_3__259_, data_stage_3__258_, data_stage_3__257_, data_stage_3__256_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__511_, data_stage_4__510_, data_stage_4__509_, data_stage_4__508_, data_stage_4__507_, data_stage_4__506_, data_stage_4__505_, data_stage_4__504_, data_stage_4__503_, data_stage_4__502_, data_stage_4__501_, data_stage_4__500_, data_stage_4__499_, data_stage_4__498_, data_stage_4__497_, data_stage_4__496_, data_stage_4__495_, data_stage_4__494_, data_stage_4__493_, data_stage_4__492_, data_stage_4__491_, data_stage_4__490_, data_stage_4__489_, data_stage_4__488_, data_stage_4__487_, data_stage_4__486_, data_stage_4__485_, data_stage_4__484_, data_stage_4__483_, data_stage_4__482_, data_stage_4__481_, data_stage_4__480_, data_stage_4__479_, data_stage_4__478_, data_stage_4__477_, data_stage_4__476_, data_stage_4__475_, data_stage_4__474_, data_stage_4__473_, data_stage_4__472_, data_stage_4__471_, data_stage_4__470_, data_stage_4__469_, data_stage_4__468_, data_stage_4__467_, data_stage_4__466_, data_stage_4__465_, data_stage_4__464_, data_stage_4__463_, data_stage_4__462_, data_stage_4__461_, data_stage_4__460_, data_stage_4__459_, data_stage_4__458_, data_stage_4__457_, data_stage_4__456_, data_stage_4__455_, data_stage_4__454_, data_stage_4__453_, data_stage_4__452_, data_stage_4__451_, data_stage_4__450_, data_stage_4__449_, data_stage_4__448_, data_stage_4__447_, data_stage_4__446_, data_stage_4__445_, data_stage_4__444_, data_stage_4__443_, data_stage_4__442_, data_stage_4__441_, data_stage_4__440_, data_stage_4__439_, data_stage_4__438_, data_stage_4__437_, data_stage_4__436_, data_stage_4__435_, data_stage_4__434_, data_stage_4__433_, data_stage_4__432_, data_stage_4__431_, data_stage_4__430_, data_stage_4__429_, data_stage_4__428_, data_stage_4__427_, data_stage_4__426_, data_stage_4__425_, data_stage_4__424_, data_stage_4__423_, data_stage_4__422_, data_stage_4__421_, data_stage_4__420_, data_stage_4__419_, data_stage_4__418_, data_stage_4__417_, data_stage_4__416_, data_stage_4__415_, data_stage_4__414_, data_stage_4__413_, data_stage_4__412_, data_stage_4__411_, data_stage_4__410_, data_stage_4__409_, data_stage_4__408_, data_stage_4__407_, data_stage_4__406_, data_stage_4__405_, data_stage_4__404_, data_stage_4__403_, data_stage_4__402_, data_stage_4__401_, data_stage_4__400_, data_stage_4__399_, data_stage_4__398_, data_stage_4__397_, data_stage_4__396_, data_stage_4__395_, data_stage_4__394_, data_stage_4__393_, data_stage_4__392_, data_stage_4__391_, data_stage_4__390_, data_stage_4__389_, data_stage_4__388_, data_stage_4__387_, data_stage_4__386_, data_stage_4__385_, data_stage_4__384_, data_stage_4__383_, data_stage_4__382_, data_stage_4__381_, data_stage_4__380_, data_stage_4__379_, data_stage_4__378_, data_stage_4__377_, data_stage_4__376_, data_stage_4__375_, data_stage_4__374_, data_stage_4__373_, data_stage_4__372_, data_stage_4__371_, data_stage_4__370_, data_stage_4__369_, data_stage_4__368_, data_stage_4__367_, data_stage_4__366_, data_stage_4__365_, data_stage_4__364_, data_stage_4__363_, data_stage_4__362_, data_stage_4__361_, data_stage_4__360_, data_stage_4__359_, data_stage_4__358_, data_stage_4__357_, data_stage_4__356_, data_stage_4__355_, data_stage_4__354_, data_stage_4__353_, data_stage_4__352_, data_stage_4__351_, data_stage_4__350_, data_stage_4__349_, data_stage_4__348_, data_stage_4__347_, data_stage_4__346_, data_stage_4__345_, data_stage_4__344_, data_stage_4__343_, data_stage_4__342_, data_stage_4__341_, data_stage_4__340_, data_stage_4__339_, data_stage_4__338_, data_stage_4__337_, data_stage_4__336_, data_stage_4__335_, data_stage_4__334_, data_stage_4__333_, data_stage_4__332_, data_stage_4__331_, data_stage_4__330_, data_stage_4__329_, data_stage_4__328_, data_stage_4__327_, data_stage_4__326_, data_stage_4__325_, data_stage_4__324_, data_stage_4__323_, data_stage_4__322_, data_stage_4__321_, data_stage_4__320_, data_stage_4__319_, data_stage_4__318_, data_stage_4__317_, data_stage_4__316_, data_stage_4__315_, data_stage_4__314_, data_stage_4__313_, data_stage_4__312_, data_stage_4__311_, data_stage_4__310_, data_stage_4__309_, data_stage_4__308_, data_stage_4__307_, data_stage_4__306_, data_stage_4__305_, data_stage_4__304_, data_stage_4__303_, data_stage_4__302_, data_stage_4__301_, data_stage_4__300_, data_stage_4__299_, data_stage_4__298_, data_stage_4__297_, data_stage_4__296_, data_stage_4__295_, data_stage_4__294_, data_stage_4__293_, data_stage_4__292_, data_stage_4__291_, data_stage_4__290_, data_stage_4__289_, data_stage_4__288_, data_stage_4__287_, data_stage_4__286_, data_stage_4__285_, data_stage_4__284_, data_stage_4__283_, data_stage_4__282_, data_stage_4__281_, data_stage_4__280_, data_stage_4__279_, data_stage_4__278_, data_stage_4__277_, data_stage_4__276_, data_stage_4__275_, data_stage_4__274_, data_stage_4__273_, data_stage_4__272_, data_stage_4__271_, data_stage_4__270_, data_stage_4__269_, data_stage_4__268_, data_stage_4__267_, data_stage_4__266_, data_stage_4__265_, data_stage_4__264_, data_stage_4__263_, data_stage_4__262_, data_stage_4__261_, data_stage_4__260_, data_stage_4__259_, data_stage_4__258_, data_stage_4__257_, data_stage_4__256_ })
  );


  bsg_swap_width_p256
  \mux_stage_4_.mux_swap_0_.swap_inst 
  (
    .data_i({ data_stage_4__511_, data_stage_4__510_, data_stage_4__509_, data_stage_4__508_, data_stage_4__507_, data_stage_4__506_, data_stage_4__505_, data_stage_4__504_, data_stage_4__503_, data_stage_4__502_, data_stage_4__501_, data_stage_4__500_, data_stage_4__499_, data_stage_4__498_, data_stage_4__497_, data_stage_4__496_, data_stage_4__495_, data_stage_4__494_, data_stage_4__493_, data_stage_4__492_, data_stage_4__491_, data_stage_4__490_, data_stage_4__489_, data_stage_4__488_, data_stage_4__487_, data_stage_4__486_, data_stage_4__485_, data_stage_4__484_, data_stage_4__483_, data_stage_4__482_, data_stage_4__481_, data_stage_4__480_, data_stage_4__479_, data_stage_4__478_, data_stage_4__477_, data_stage_4__476_, data_stage_4__475_, data_stage_4__474_, data_stage_4__473_, data_stage_4__472_, data_stage_4__471_, data_stage_4__470_, data_stage_4__469_, data_stage_4__468_, data_stage_4__467_, data_stage_4__466_, data_stage_4__465_, data_stage_4__464_, data_stage_4__463_, data_stage_4__462_, data_stage_4__461_, data_stage_4__460_, data_stage_4__459_, data_stage_4__458_, data_stage_4__457_, data_stage_4__456_, data_stage_4__455_, data_stage_4__454_, data_stage_4__453_, data_stage_4__452_, data_stage_4__451_, data_stage_4__450_, data_stage_4__449_, data_stage_4__448_, data_stage_4__447_, data_stage_4__446_, data_stage_4__445_, data_stage_4__444_, data_stage_4__443_, data_stage_4__442_, data_stage_4__441_, data_stage_4__440_, data_stage_4__439_, data_stage_4__438_, data_stage_4__437_, data_stage_4__436_, data_stage_4__435_, data_stage_4__434_, data_stage_4__433_, data_stage_4__432_, data_stage_4__431_, data_stage_4__430_, data_stage_4__429_, data_stage_4__428_, data_stage_4__427_, data_stage_4__426_, data_stage_4__425_, data_stage_4__424_, data_stage_4__423_, data_stage_4__422_, data_stage_4__421_, data_stage_4__420_, data_stage_4__419_, data_stage_4__418_, data_stage_4__417_, data_stage_4__416_, data_stage_4__415_, data_stage_4__414_, data_stage_4__413_, data_stage_4__412_, data_stage_4__411_, data_stage_4__410_, data_stage_4__409_, data_stage_4__408_, data_stage_4__407_, data_stage_4__406_, data_stage_4__405_, data_stage_4__404_, data_stage_4__403_, data_stage_4__402_, data_stage_4__401_, data_stage_4__400_, data_stage_4__399_, data_stage_4__398_, data_stage_4__397_, data_stage_4__396_, data_stage_4__395_, data_stage_4__394_, data_stage_4__393_, data_stage_4__392_, data_stage_4__391_, data_stage_4__390_, data_stage_4__389_, data_stage_4__388_, data_stage_4__387_, data_stage_4__386_, data_stage_4__385_, data_stage_4__384_, data_stage_4__383_, data_stage_4__382_, data_stage_4__381_, data_stage_4__380_, data_stage_4__379_, data_stage_4__378_, data_stage_4__377_, data_stage_4__376_, data_stage_4__375_, data_stage_4__374_, data_stage_4__373_, data_stage_4__372_, data_stage_4__371_, data_stage_4__370_, data_stage_4__369_, data_stage_4__368_, data_stage_4__367_, data_stage_4__366_, data_stage_4__365_, data_stage_4__364_, data_stage_4__363_, data_stage_4__362_, data_stage_4__361_, data_stage_4__360_, data_stage_4__359_, data_stage_4__358_, data_stage_4__357_, data_stage_4__356_, data_stage_4__355_, data_stage_4__354_, data_stage_4__353_, data_stage_4__352_, data_stage_4__351_, data_stage_4__350_, data_stage_4__349_, data_stage_4__348_, data_stage_4__347_, data_stage_4__346_, data_stage_4__345_, data_stage_4__344_, data_stage_4__343_, data_stage_4__342_, data_stage_4__341_, data_stage_4__340_, data_stage_4__339_, data_stage_4__338_, data_stage_4__337_, data_stage_4__336_, data_stage_4__335_, data_stage_4__334_, data_stage_4__333_, data_stage_4__332_, data_stage_4__331_, data_stage_4__330_, data_stage_4__329_, data_stage_4__328_, data_stage_4__327_, data_stage_4__326_, data_stage_4__325_, data_stage_4__324_, data_stage_4__323_, data_stage_4__322_, data_stage_4__321_, data_stage_4__320_, data_stage_4__319_, data_stage_4__318_, data_stage_4__317_, data_stage_4__316_, data_stage_4__315_, data_stage_4__314_, data_stage_4__313_, data_stage_4__312_, data_stage_4__311_, data_stage_4__310_, data_stage_4__309_, data_stage_4__308_, data_stage_4__307_, data_stage_4__306_, data_stage_4__305_, data_stage_4__304_, data_stage_4__303_, data_stage_4__302_, data_stage_4__301_, data_stage_4__300_, data_stage_4__299_, data_stage_4__298_, data_stage_4__297_, data_stage_4__296_, data_stage_4__295_, data_stage_4__294_, data_stage_4__293_, data_stage_4__292_, data_stage_4__291_, data_stage_4__290_, data_stage_4__289_, data_stage_4__288_, data_stage_4__287_, data_stage_4__286_, data_stage_4__285_, data_stage_4__284_, data_stage_4__283_, data_stage_4__282_, data_stage_4__281_, data_stage_4__280_, data_stage_4__279_, data_stage_4__278_, data_stage_4__277_, data_stage_4__276_, data_stage_4__275_, data_stage_4__274_, data_stage_4__273_, data_stage_4__272_, data_stage_4__271_, data_stage_4__270_, data_stage_4__269_, data_stage_4__268_, data_stage_4__267_, data_stage_4__266_, data_stage_4__265_, data_stage_4__264_, data_stage_4__263_, data_stage_4__262_, data_stage_4__261_, data_stage_4__260_, data_stage_4__259_, data_stage_4__258_, data_stage_4__257_, data_stage_4__256_, data_stage_4__255_, data_stage_4__254_, data_stage_4__253_, data_stage_4__252_, data_stage_4__251_, data_stage_4__250_, data_stage_4__249_, data_stage_4__248_, data_stage_4__247_, data_stage_4__246_, data_stage_4__245_, data_stage_4__244_, data_stage_4__243_, data_stage_4__242_, data_stage_4__241_, data_stage_4__240_, data_stage_4__239_, data_stage_4__238_, data_stage_4__237_, data_stage_4__236_, data_stage_4__235_, data_stage_4__234_, data_stage_4__233_, data_stage_4__232_, data_stage_4__231_, data_stage_4__230_, data_stage_4__229_, data_stage_4__228_, data_stage_4__227_, data_stage_4__226_, data_stage_4__225_, data_stage_4__224_, data_stage_4__223_, data_stage_4__222_, data_stage_4__221_, data_stage_4__220_, data_stage_4__219_, data_stage_4__218_, data_stage_4__217_, data_stage_4__216_, data_stage_4__215_, data_stage_4__214_, data_stage_4__213_, data_stage_4__212_, data_stage_4__211_, data_stage_4__210_, data_stage_4__209_, data_stage_4__208_, data_stage_4__207_, data_stage_4__206_, data_stage_4__205_, data_stage_4__204_, data_stage_4__203_, data_stage_4__202_, data_stage_4__201_, data_stage_4__200_, data_stage_4__199_, data_stage_4__198_, data_stage_4__197_, data_stage_4__196_, data_stage_4__195_, data_stage_4__194_, data_stage_4__193_, data_stage_4__192_, data_stage_4__191_, data_stage_4__190_, data_stage_4__189_, data_stage_4__188_, data_stage_4__187_, data_stage_4__186_, data_stage_4__185_, data_stage_4__184_, data_stage_4__183_, data_stage_4__182_, data_stage_4__181_, data_stage_4__180_, data_stage_4__179_, data_stage_4__178_, data_stage_4__177_, data_stage_4__176_, data_stage_4__175_, data_stage_4__174_, data_stage_4__173_, data_stage_4__172_, data_stage_4__171_, data_stage_4__170_, data_stage_4__169_, data_stage_4__168_, data_stage_4__167_, data_stage_4__166_, data_stage_4__165_, data_stage_4__164_, data_stage_4__163_, data_stage_4__162_, data_stage_4__161_, data_stage_4__160_, data_stage_4__159_, data_stage_4__158_, data_stage_4__157_, data_stage_4__156_, data_stage_4__155_, data_stage_4__154_, data_stage_4__153_, data_stage_4__152_, data_stage_4__151_, data_stage_4__150_, data_stage_4__149_, data_stage_4__148_, data_stage_4__147_, data_stage_4__146_, data_stage_4__145_, data_stage_4__144_, data_stage_4__143_, data_stage_4__142_, data_stage_4__141_, data_stage_4__140_, data_stage_4__139_, data_stage_4__138_, data_stage_4__137_, data_stage_4__136_, data_stage_4__135_, data_stage_4__134_, data_stage_4__133_, data_stage_4__132_, data_stage_4__131_, data_stage_4__130_, data_stage_4__129_, data_stage_4__128_, data_stage_4__127_, data_stage_4__126_, data_stage_4__125_, data_stage_4__124_, data_stage_4__123_, data_stage_4__122_, data_stage_4__121_, data_stage_4__120_, data_stage_4__119_, data_stage_4__118_, data_stage_4__117_, data_stage_4__116_, data_stage_4__115_, data_stage_4__114_, data_stage_4__113_, data_stage_4__112_, data_stage_4__111_, data_stage_4__110_, data_stage_4__109_, data_stage_4__108_, data_stage_4__107_, data_stage_4__106_, data_stage_4__105_, data_stage_4__104_, data_stage_4__103_, data_stage_4__102_, data_stage_4__101_, data_stage_4__100_, data_stage_4__99_, data_stage_4__98_, data_stage_4__97_, data_stage_4__96_, data_stage_4__95_, data_stage_4__94_, data_stage_4__93_, data_stage_4__92_, data_stage_4__91_, data_stage_4__90_, data_stage_4__89_, data_stage_4__88_, data_stage_4__87_, data_stage_4__86_, data_stage_4__85_, data_stage_4__84_, data_stage_4__83_, data_stage_4__82_, data_stage_4__81_, data_stage_4__80_, data_stage_4__79_, data_stage_4__78_, data_stage_4__77_, data_stage_4__76_, data_stage_4__75_, data_stage_4__74_, data_stage_4__73_, data_stage_4__72_, data_stage_4__71_, data_stage_4__70_, data_stage_4__69_, data_stage_4__68_, data_stage_4__67_, data_stage_4__66_, data_stage_4__65_, data_stage_4__64_, data_stage_4__63_, data_stage_4__62_, data_stage_4__61_, data_stage_4__60_, data_stage_4__59_, data_stage_4__58_, data_stage_4__57_, data_stage_4__56_, data_stage_4__55_, data_stage_4__54_, data_stage_4__53_, data_stage_4__52_, data_stage_4__51_, data_stage_4__50_, data_stage_4__49_, data_stage_4__48_, data_stage_4__47_, data_stage_4__46_, data_stage_4__45_, data_stage_4__44_, data_stage_4__43_, data_stage_4__42_, data_stage_4__41_, data_stage_4__40_, data_stage_4__39_, data_stage_4__38_, data_stage_4__37_, data_stage_4__36_, data_stage_4__35_, data_stage_4__34_, data_stage_4__33_, data_stage_4__32_, data_stage_4__31_, data_stage_4__30_, data_stage_4__29_, data_stage_4__28_, data_stage_4__27_, data_stage_4__26_, data_stage_4__25_, data_stage_4__24_, data_stage_4__23_, data_stage_4__22_, data_stage_4__21_, data_stage_4__20_, data_stage_4__19_, data_stage_4__18_, data_stage_4__17_, data_stage_4__16_, data_stage_4__15_, data_stage_4__14_, data_stage_4__13_, data_stage_4__12_, data_stage_4__11_, data_stage_4__10_, data_stage_4__9_, data_stage_4__8_, data_stage_4__7_, data_stage_4__6_, data_stage_4__5_, data_stage_4__4_, data_stage_4__3_, data_stage_4__2_, data_stage_4__1_, data_stage_4__0_ }),
    .swap_i(sel_i[4]),
    .data_o(data_o)
  );


endmodule

